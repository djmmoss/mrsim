module Fifo_0(input clk, input reset,
    input  io_enq_val,
    output io_enq_rdy,
    output io_deq_val,
    input  io_deq_rdy,
    input [63:0] io_enq_dat,
    output[63:0] io_deq_dat
);

  wire[63:0] T0;
  wire[63:0] T1;
  reg [63:0] ram [3:0];
  wire[63:0] T2;
  wire[63:0] T3;
  wire do_enq;
  wire T4;
  reg[0:0] is_full;
  wire is_full_next;
  wire T5;
  wire T6;
  wire do_deq;
  wire T7;
  wire is_empty;
  wire T8;
  reg[3:0] deq_ptr;
  wire[3:0] T9;
  wire[3:0] deq_ptr_inc;
  reg[3:0] enq_ptr;
  wire[3:0] T10;
  wire[3:0] enq_ptr_inc;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;

  assign io_deq_dat = T0;
  assign T0 = do_deq ? T1 : 64'h0;
  assign T1 = ram[T17];
  assign T3 = io_enq_dat;
  assign do_enq = T4 && io_enq_val;
  assign T4 = ! is_full;
  assign is_full_next = T12 ? 1'h1 : T5;
  assign T5 = T6 ? 1'h0 : is_full;
  assign T6 = do_deq && is_full;
  assign do_deq = io_deq_rdy && T7;
  assign T7 = ! is_empty;
  assign is_empty = T11 && T8;
  assign T8 = enq_ptr == deq_ptr;
  assign T9 = do_deq ? deq_ptr_inc : deq_ptr;
  assign deq_ptr_inc = deq_ptr + 4'h1;
  assign T10 = do_enq ? enq_ptr_inc : enq_ptr;
  assign enq_ptr_inc = enq_ptr + 4'h1;
  assign T11 = ! is_full;
  assign T12 = T14 && T13;
  assign T13 = enq_ptr_inc == deq_ptr;
  assign T14 = do_enq && T15;
  assign T15 = ~ do_deq;
  assign T16 = enq_ptr[1'h1:1'h0];
  assign T17 = deq_ptr[1'h1:1'h0];
  assign io_deq_val = T18;
  assign T18 = ! is_empty;
  assign io_enq_rdy = T19;
  assign T19 = ! is_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[T16] <= T3;
    is_full <= reset ? 1'h0 : is_full_next;
    deq_ptr <= reset ? 4'h0 : T9;
    enq_ptr <= reset ? 4'h0 : T10;
  end
endmodule

module encode(
    input [63:0] io_rx_dat_int,
    output io_rx_rdy,
    input  io_rx_val,
    output[63:0] io_tx_dat,
    output io_tx_val
);


  assign io_tx_val = io_rx_val;
  assign io_tx_dat = io_rx_dat_int;
  assign io_rx_rdy = 1'h1;
endmodule

module decode(
    input [63:0] io_rx_dat,
    output io_rx_rdy,
    input  io_rx_val,
    output[63:0] io_tx_dat_int,
    output io_tx_val
);


  assign io_tx_val = io_rx_val;
  assign io_tx_dat_int = io_rx_dat;
  assign io_rx_rdy = 1'h1;
endmodule

module Fifo_1(input clk, input reset,
    input  io_enq_val,
    output io_enq_rdy,
    output io_deq_val,
    input  io_deq_rdy,
    input [63:0] io_enq_dat_int,
    output[63:0] io_deq_dat_int
);

  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [63:0] ram [3:0];
  wire[63:0] T4;
  wire[63:0] T5;
  wire do_enq;
  wire T6;
  reg[0:0] is_full;
  wire is_full_next;
  wire T7;
  wire T8;
  wire do_deq;
  wire T9;
  wire is_empty;
  wire T10;
  reg[3:0] deq_ptr;
  wire[3:0] T11;
  wire[3:0] deq_ptr_inc;
  reg[3:0] enq_ptr;
  wire[3:0] T12;
  wire[3:0] enq_ptr_inc;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;

  assign io_deq_dat_int = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = do_deq ? T2 : 64'h0;
  assign T2 = T3[6'h3f:1'h0];
  assign T3 = ram[T19];
  assign T5 = io_enq_dat_int;
  assign do_enq = T6 && io_enq_val;
  assign T6 = ! is_full;
  assign is_full_next = T14 ? 1'h1 : T7;
  assign T7 = T8 ? 1'h0 : is_full;
  assign T8 = do_deq && is_full;
  assign do_deq = io_deq_rdy && T9;
  assign T9 = ! is_empty;
  assign is_empty = T13 && T10;
  assign T10 = enq_ptr == deq_ptr;
  assign T11 = do_deq ? deq_ptr_inc : deq_ptr;
  assign deq_ptr_inc = deq_ptr + 4'h1;
  assign T12 = do_enq ? enq_ptr_inc : enq_ptr;
  assign enq_ptr_inc = enq_ptr + 4'h1;
  assign T13 = ! is_full;
  assign T14 = T16 && T15;
  assign T15 = enq_ptr_inc == deq_ptr;
  assign T16 = do_enq && T17;
  assign T17 = ~ do_deq;
  assign T18 = enq_ptr[1'h1:1'h0];
  assign T19 = deq_ptr[1'h1:1'h0];
  assign io_deq_val = T20;
  assign T20 = ! is_empty;
  assign io_enq_rdy = T21;
  assign T21 = ! is_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[T18] <= T5;
    is_full <= reset ? 1'h0 : is_full_next;
    deq_ptr <= reset ? 4'h0 : T11;
    enq_ptr <= reset ? 4'h0 : T12;
  end
endmodule

module Cell(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;

  assign io_out = isAlive;
  assign T0 = T40 || T1;
  assign T1 = T39 && T2;
  assign T2 = T30 && T3;
  assign T3 = T29 && T4;
  assign T4 = count == 3'h3;
  assign count = T27 + T5;
  assign T5 = T25 + T6;
  assign T6 = T23 + T7;
  assign T7 = T21 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T19 + T10;
  assign T10 = T17 + T11;
  assign T11 = T15 + T12;
  assign T12 = T13 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_8;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_7;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_6;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_5;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_3;
  assign T23 = {2'h0, T24};
  assign T24 = io_nbrs_2;
  assign T25 = {2'h0, T26};
  assign T26 = io_nbrs_1;
  assign T27 = {2'h0, T28};
  assign T28 = io_nbrs_0;
  assign T29 = ! isAlive;
  assign T30 = ! T31;
  assign T31 = T34 || T32;
  assign T32 = isAlive && T33;
  assign T33 = 3'h4 <= count;
  assign T34 = T37 || T35;
  assign T35 = isAlive && T36;
  assign T36 = count < 3'h4;
  assign T37 = isAlive && T38;
  assign T38 = count < 3'h2;
  assign T39 = ! io_in_val;
  assign T40 = T44 || T41;
  assign T41 = T39 && T42;
  assign T42 = T43 && T32;
  assign T43 = ! T34;
  assign T44 = T48 || T45;
  assign T45 = T39 && T46;
  assign T46 = T47 && T35;
  assign T47 = ! T37;
  assign T48 = io_in_val || T49;
  assign T49 = T39 && T37;
  assign T50 = T1 ? 1'h1 : T51;
  assign T51 = T41 ? 1'h0 : T52;
  assign T52 = T45 ? 1'h1 : T53;
  assign T53 = T49 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T50;
    end
  end
endmodule

module Mapper(input clk, input reset,
    input [63:0] io_rx_dat_int,
    input  io_rx_val,
    output io_rx_rdy,
    output[63:0] io_tx_dat_int,
    output io_tx_val
);

  wire Cell_0_io_out;
  wire Cell_7_io_out;
  wire Cell_6_io_out;
  wire Cell_56_io_out;
  wire Cell_62_io_out;
  wire Cell_48_io_out;
  wire Cell_55_io_out;
  wire Cell_54_io_out;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[63:0] in;
  wire Cell_63_io_out;
  wire Cell_40_io_out;
  wire Cell_47_io_out;
  wire Cell_46_io_out;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire Cell_32_io_out;
  wire Cell_39_io_out;
  wire Cell_38_io_out;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire Cell_24_io_out;
  wire Cell_31_io_out;
  wire Cell_30_io_out;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire Cell_16_io_out;
  wire Cell_23_io_out;
  wire Cell_22_io_out;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire Cell_8_io_out;
  wire Cell_15_io_out;
  wire Cell_14_io_out;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire Cell_5_io_out;
  wire Cell_61_io_out;
  wire Cell_53_io_out;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire Cell_45_io_out;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire Cell_37_io_out;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire Cell_29_io_out;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire Cell_21_io_out;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire Cell_13_io_out;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire Cell_4_io_out;
  wire Cell_60_io_out;
  wire Cell_52_io_out;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire Cell_44_io_out;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire Cell_36_io_out;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire Cell_28_io_out;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire Cell_20_io_out;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire Cell_12_io_out;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire Cell_3_io_out;
  wire Cell_59_io_out;
  wire Cell_51_io_out;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire Cell_43_io_out;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire Cell_35_io_out;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire Cell_27_io_out;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire Cell_19_io_out;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire Cell_11_io_out;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire Cell_2_io_out;
  wire Cell_58_io_out;
  wire Cell_50_io_out;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire Cell_42_io_out;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire Cell_34_io_out;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire Cell_26_io_out;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire Cell_18_io_out;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire Cell_10_io_out;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire Cell_1_io_out;
  wire Cell_57_io_out;
  wire Cell_49_io_out;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire Cell_41_io_out;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire Cell_33_io_out;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire Cell_25_io_out;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire Cell_17_io_out;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire Cell_9_io_out;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  reg[6:0] R386;
  wire[6:0] T387;
  wire[6:0] T388;
  wire T389;
  wire T390;
  wire[63:0] T391;
  wire[63:0] T392;
  reg[63:0] check_out;
  wire T393;
  wire[63:0] T394;
  wire[63:0] T395;
  wire[63:0] T396;
  wire[63:0] T397;
  wire out_0;
  wire[62:0] T398;
  wire out_1;
  wire[61:0] T399;
  wire out_2;
  wire[60:0] T400;
  wire out_3;
  wire[59:0] T401;
  wire out_4;
  wire[58:0] T402;
  wire out_5;
  wire[57:0] T403;
  wire out_6;
  wire[56:0] T404;
  wire out_7;
  wire[55:0] T405;
  wire out_8;
  wire[54:0] T406;
  wire out_9;
  wire[53:0] T407;
  wire out_10;
  wire[52:0] T408;
  wire out_11;
  wire[51:0] T409;
  wire out_12;
  wire[50:0] T410;
  wire out_13;
  wire[49:0] T411;
  wire out_14;
  wire[48:0] T412;
  wire out_15;
  wire[47:0] T413;
  wire out_16;
  wire[46:0] T414;
  wire out_17;
  wire[45:0] T415;
  wire out_18;
  wire[44:0] T416;
  wire out_19;
  wire[43:0] T417;
  wire out_20;
  wire[42:0] T418;
  wire out_21;
  wire[41:0] T419;
  wire out_22;
  wire[40:0] T420;
  wire out_23;
  wire[39:0] T421;
  wire out_24;
  wire[38:0] T422;
  wire out_25;
  wire[37:0] T423;
  wire out_26;
  wire[36:0] T424;
  wire out_27;
  wire[35:0] T425;
  wire out_28;
  wire[34:0] T426;
  wire out_29;
  wire[33:0] T427;
  wire out_30;
  wire[32:0] T428;
  wire out_31;
  wire[31:0] T429;
  wire out_32;
  wire[30:0] T430;
  wire out_33;
  wire[29:0] T431;
  wire out_34;
  wire[28:0] T432;
  wire out_35;
  wire[27:0] T433;
  wire out_36;
  wire[26:0] T434;
  wire out_37;
  wire[25:0] T435;
  wire out_38;
  wire[24:0] T436;
  wire out_39;
  wire[23:0] T437;
  wire out_40;
  wire[22:0] T438;
  wire out_41;
  wire[21:0] T439;
  wire out_42;
  wire[20:0] T440;
  wire out_43;
  wire[19:0] T441;
  wire out_44;
  wire[18:0] T442;
  wire out_45;
  wire[17:0] T443;
  wire out_46;
  wire[16:0] T444;
  wire out_47;
  wire[15:0] T445;
  wire out_48;
  wire[14:0] T446;
  wire out_49;
  wire[13:0] T447;
  wire out_50;
  wire[12:0] T448;
  wire out_51;
  wire[11:0] T449;
  wire out_52;
  wire[10:0] T450;
  wire out_53;
  wire[9:0] T451;
  wire out_54;
  wire[8:0] T452;
  wire out_55;
  wire[7:0] T453;
  wire out_56;
  wire[6:0] T454;
  wire out_57;
  wire[5:0] T455;
  wire out_58;
  wire[4:0] T456;
  wire out_59;
  wire[3:0] T457;
  wire out_60;
  wire[2:0] T458;
  wire out_61;
  wire[1:0] T459;
  wire out_62;
  wire out_63;
  wire T460;
  reg[0:0] is_full;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;

  assign T0 = T1 ? 1'h0 : io_rx_val;
  assign T1 = ! io_rx_val;
  assign T2 = T1 ? 1'h0 : T3;
  assign T3 = io_rx_val ? T4 : 1'h0;
  assign T4 = T5;
  assign T5 = in[6'h3f:6'h3f];
  assign in = io_rx_dat_int;
  assign T6 = T7 ? 1'h0 : io_rx_val;
  assign T7 = ! io_rx_val;
  assign T8 = T7 ? 1'h0 : T9;
  assign T9 = io_rx_val ? T10 : 1'h0;
  assign T10 = T11;
  assign T11 = in[6'h3e:6'h3e];
  assign T12 = T13 ? 1'h0 : io_rx_val;
  assign T13 = ! io_rx_val;
  assign T14 = T13 ? 1'h0 : T15;
  assign T15 = io_rx_val ? T16 : 1'h0;
  assign T16 = T17;
  assign T17 = in[6'h3d:6'h3d];
  assign T18 = T19 ? 1'h0 : io_rx_val;
  assign T19 = ! io_rx_val;
  assign T20 = T19 ? 1'h0 : T21;
  assign T21 = io_rx_val ? T22 : 1'h0;
  assign T22 = T23;
  assign T23 = in[6'h3c:6'h3c];
  assign T24 = T25 ? 1'h0 : io_rx_val;
  assign T25 = ! io_rx_val;
  assign T26 = T25 ? 1'h0 : T27;
  assign T27 = io_rx_val ? T28 : 1'h0;
  assign T28 = T29;
  assign T29 = in[6'h3b:6'h3b];
  assign T30 = T31 ? 1'h0 : io_rx_val;
  assign T31 = ! io_rx_val;
  assign T32 = T31 ? 1'h0 : T33;
  assign T33 = io_rx_val ? T34 : 1'h0;
  assign T34 = T35;
  assign T35 = in[6'h3a:6'h3a];
  assign T36 = T37 ? 1'h0 : io_rx_val;
  assign T37 = ! io_rx_val;
  assign T38 = T37 ? 1'h0 : T39;
  assign T39 = io_rx_val ? T40 : 1'h0;
  assign T40 = T41;
  assign T41 = in[6'h39:6'h39];
  assign T42 = T43 ? 1'h0 : io_rx_val;
  assign T43 = ! io_rx_val;
  assign T44 = T43 ? 1'h0 : T45;
  assign T45 = io_rx_val ? T46 : 1'h0;
  assign T46 = T47;
  assign T47 = in[6'h38:6'h38];
  assign T48 = T49 ? 1'h0 : io_rx_val;
  assign T49 = ! io_rx_val;
  assign T50 = T49 ? 1'h0 : T51;
  assign T51 = io_rx_val ? T52 : 1'h0;
  assign T52 = T53;
  assign T53 = in[6'h37:6'h37];
  assign T54 = T55 ? 1'h0 : io_rx_val;
  assign T55 = ! io_rx_val;
  assign T56 = T55 ? 1'h0 : T57;
  assign T57 = io_rx_val ? T58 : 1'h0;
  assign T58 = T59;
  assign T59 = in[6'h36:6'h36];
  assign T60 = T61 ? 1'h0 : io_rx_val;
  assign T61 = ! io_rx_val;
  assign T62 = T61 ? 1'h0 : T63;
  assign T63 = io_rx_val ? T64 : 1'h0;
  assign T64 = T65;
  assign T65 = in[6'h35:6'h35];
  assign T66 = T67 ? 1'h0 : io_rx_val;
  assign T67 = ! io_rx_val;
  assign T68 = T67 ? 1'h0 : T69;
  assign T69 = io_rx_val ? T70 : 1'h0;
  assign T70 = T71;
  assign T71 = in[6'h34:6'h34];
  assign T72 = T73 ? 1'h0 : io_rx_val;
  assign T73 = ! io_rx_val;
  assign T74 = T73 ? 1'h0 : T75;
  assign T75 = io_rx_val ? T76 : 1'h0;
  assign T76 = T77;
  assign T77 = in[6'h33:6'h33];
  assign T78 = T79 ? 1'h0 : io_rx_val;
  assign T79 = ! io_rx_val;
  assign T80 = T79 ? 1'h0 : T81;
  assign T81 = io_rx_val ? T82 : 1'h0;
  assign T82 = T83;
  assign T83 = in[6'h32:6'h32];
  assign T84 = T85 ? 1'h0 : io_rx_val;
  assign T85 = ! io_rx_val;
  assign T86 = T85 ? 1'h0 : T87;
  assign T87 = io_rx_val ? T88 : 1'h0;
  assign T88 = T89;
  assign T89 = in[6'h31:6'h31];
  assign T90 = T91 ? 1'h0 : io_rx_val;
  assign T91 = ! io_rx_val;
  assign T92 = T91 ? 1'h0 : T93;
  assign T93 = io_rx_val ? T94 : 1'h0;
  assign T94 = T95;
  assign T95 = in[6'h30:6'h30];
  assign T96 = T97 ? 1'h0 : io_rx_val;
  assign T97 = ! io_rx_val;
  assign T98 = T97 ? 1'h0 : T99;
  assign T99 = io_rx_val ? T100 : 1'h0;
  assign T100 = T101;
  assign T101 = in[6'h2f:6'h2f];
  assign T102 = T103 ? 1'h0 : io_rx_val;
  assign T103 = ! io_rx_val;
  assign T104 = T103 ? 1'h0 : T105;
  assign T105 = io_rx_val ? T106 : 1'h0;
  assign T106 = T107;
  assign T107 = in[6'h2e:6'h2e];
  assign T108 = T109 ? 1'h0 : io_rx_val;
  assign T109 = ! io_rx_val;
  assign T110 = T109 ? 1'h0 : T111;
  assign T111 = io_rx_val ? T112 : 1'h0;
  assign T112 = T113;
  assign T113 = in[6'h2d:6'h2d];
  assign T114 = T115 ? 1'h0 : io_rx_val;
  assign T115 = ! io_rx_val;
  assign T116 = T115 ? 1'h0 : T117;
  assign T117 = io_rx_val ? T118 : 1'h0;
  assign T118 = T119;
  assign T119 = in[6'h2c:6'h2c];
  assign T120 = T121 ? 1'h0 : io_rx_val;
  assign T121 = ! io_rx_val;
  assign T122 = T121 ? 1'h0 : T123;
  assign T123 = io_rx_val ? T124 : 1'h0;
  assign T124 = T125;
  assign T125 = in[6'h2b:6'h2b];
  assign T126 = T127 ? 1'h0 : io_rx_val;
  assign T127 = ! io_rx_val;
  assign T128 = T127 ? 1'h0 : T129;
  assign T129 = io_rx_val ? T130 : 1'h0;
  assign T130 = T131;
  assign T131 = in[6'h2a:6'h2a];
  assign T132 = T133 ? 1'h0 : io_rx_val;
  assign T133 = ! io_rx_val;
  assign T134 = T133 ? 1'h0 : T135;
  assign T135 = io_rx_val ? T136 : 1'h0;
  assign T136 = T137;
  assign T137 = in[6'h29:6'h29];
  assign T138 = T139 ? 1'h0 : io_rx_val;
  assign T139 = ! io_rx_val;
  assign T140 = T139 ? 1'h0 : T141;
  assign T141 = io_rx_val ? T142 : 1'h0;
  assign T142 = T143;
  assign T143 = in[6'h28:6'h28];
  assign T144 = T145 ? 1'h0 : io_rx_val;
  assign T145 = ! io_rx_val;
  assign T146 = T145 ? 1'h0 : T147;
  assign T147 = io_rx_val ? T148 : 1'h0;
  assign T148 = T149;
  assign T149 = in[6'h27:6'h27];
  assign T150 = T151 ? 1'h0 : io_rx_val;
  assign T151 = ! io_rx_val;
  assign T152 = T151 ? 1'h0 : T153;
  assign T153 = io_rx_val ? T154 : 1'h0;
  assign T154 = T155;
  assign T155 = in[6'h26:6'h26];
  assign T156 = T157 ? 1'h0 : io_rx_val;
  assign T157 = ! io_rx_val;
  assign T158 = T157 ? 1'h0 : T159;
  assign T159 = io_rx_val ? T160 : 1'h0;
  assign T160 = T161;
  assign T161 = in[6'h25:6'h25];
  assign T162 = T163 ? 1'h0 : io_rx_val;
  assign T163 = ! io_rx_val;
  assign T164 = T163 ? 1'h0 : T165;
  assign T165 = io_rx_val ? T166 : 1'h0;
  assign T166 = T167;
  assign T167 = in[6'h24:6'h24];
  assign T168 = T169 ? 1'h0 : io_rx_val;
  assign T169 = ! io_rx_val;
  assign T170 = T169 ? 1'h0 : T171;
  assign T171 = io_rx_val ? T172 : 1'h0;
  assign T172 = T173;
  assign T173 = in[6'h23:6'h23];
  assign T174 = T175 ? 1'h0 : io_rx_val;
  assign T175 = ! io_rx_val;
  assign T176 = T175 ? 1'h0 : T177;
  assign T177 = io_rx_val ? T178 : 1'h0;
  assign T178 = T179;
  assign T179 = in[6'h22:6'h22];
  assign T180 = T181 ? 1'h0 : io_rx_val;
  assign T181 = ! io_rx_val;
  assign T182 = T181 ? 1'h0 : T183;
  assign T183 = io_rx_val ? T184 : 1'h0;
  assign T184 = T185;
  assign T185 = in[6'h21:6'h21];
  assign T186 = T187 ? 1'h0 : io_rx_val;
  assign T187 = ! io_rx_val;
  assign T188 = T187 ? 1'h0 : T189;
  assign T189 = io_rx_val ? T190 : 1'h0;
  assign T190 = T191;
  assign T191 = in[6'h20:6'h20];
  assign T192 = T193 ? 1'h0 : io_rx_val;
  assign T193 = ! io_rx_val;
  assign T194 = T193 ? 1'h0 : T195;
  assign T195 = io_rx_val ? T196 : 1'h0;
  assign T196 = T197;
  assign T197 = in[5'h1f:5'h1f];
  assign T198 = T199 ? 1'h0 : io_rx_val;
  assign T199 = ! io_rx_val;
  assign T200 = T199 ? 1'h0 : T201;
  assign T201 = io_rx_val ? T202 : 1'h0;
  assign T202 = T203;
  assign T203 = in[5'h1e:5'h1e];
  assign T204 = T205 ? 1'h0 : io_rx_val;
  assign T205 = ! io_rx_val;
  assign T206 = T205 ? 1'h0 : T207;
  assign T207 = io_rx_val ? T208 : 1'h0;
  assign T208 = T209;
  assign T209 = in[5'h1d:5'h1d];
  assign T210 = T211 ? 1'h0 : io_rx_val;
  assign T211 = ! io_rx_val;
  assign T212 = T211 ? 1'h0 : T213;
  assign T213 = io_rx_val ? T214 : 1'h0;
  assign T214 = T215;
  assign T215 = in[5'h1c:5'h1c];
  assign T216 = T217 ? 1'h0 : io_rx_val;
  assign T217 = ! io_rx_val;
  assign T218 = T217 ? 1'h0 : T219;
  assign T219 = io_rx_val ? T220 : 1'h0;
  assign T220 = T221;
  assign T221 = in[5'h1b:5'h1b];
  assign T222 = T223 ? 1'h0 : io_rx_val;
  assign T223 = ! io_rx_val;
  assign T224 = T223 ? 1'h0 : T225;
  assign T225 = io_rx_val ? T226 : 1'h0;
  assign T226 = T227;
  assign T227 = in[5'h1a:5'h1a];
  assign T228 = T229 ? 1'h0 : io_rx_val;
  assign T229 = ! io_rx_val;
  assign T230 = T229 ? 1'h0 : T231;
  assign T231 = io_rx_val ? T232 : 1'h0;
  assign T232 = T233;
  assign T233 = in[5'h19:5'h19];
  assign T234 = T235 ? 1'h0 : io_rx_val;
  assign T235 = ! io_rx_val;
  assign T236 = T235 ? 1'h0 : T237;
  assign T237 = io_rx_val ? T238 : 1'h0;
  assign T238 = T239;
  assign T239 = in[5'h18:5'h18];
  assign T240 = T241 ? 1'h0 : io_rx_val;
  assign T241 = ! io_rx_val;
  assign T242 = T241 ? 1'h0 : T243;
  assign T243 = io_rx_val ? T244 : 1'h0;
  assign T244 = T245;
  assign T245 = in[5'h17:5'h17];
  assign T246 = T247 ? 1'h0 : io_rx_val;
  assign T247 = ! io_rx_val;
  assign T248 = T247 ? 1'h0 : T249;
  assign T249 = io_rx_val ? T250 : 1'h0;
  assign T250 = T251;
  assign T251 = in[5'h16:5'h16];
  assign T252 = T253 ? 1'h0 : io_rx_val;
  assign T253 = ! io_rx_val;
  assign T254 = T253 ? 1'h0 : T255;
  assign T255 = io_rx_val ? T256 : 1'h0;
  assign T256 = T257;
  assign T257 = in[5'h15:5'h15];
  assign T258 = T259 ? 1'h0 : io_rx_val;
  assign T259 = ! io_rx_val;
  assign T260 = T259 ? 1'h0 : T261;
  assign T261 = io_rx_val ? T262 : 1'h0;
  assign T262 = T263;
  assign T263 = in[5'h14:5'h14];
  assign T264 = T265 ? 1'h0 : io_rx_val;
  assign T265 = ! io_rx_val;
  assign T266 = T265 ? 1'h0 : T267;
  assign T267 = io_rx_val ? T268 : 1'h0;
  assign T268 = T269;
  assign T269 = in[5'h13:5'h13];
  assign T270 = T271 ? 1'h0 : io_rx_val;
  assign T271 = ! io_rx_val;
  assign T272 = T271 ? 1'h0 : T273;
  assign T273 = io_rx_val ? T274 : 1'h0;
  assign T274 = T275;
  assign T275 = in[5'h12:5'h12];
  assign T276 = T277 ? 1'h0 : io_rx_val;
  assign T277 = ! io_rx_val;
  assign T278 = T277 ? 1'h0 : T279;
  assign T279 = io_rx_val ? T280 : 1'h0;
  assign T280 = T281;
  assign T281 = in[5'h11:5'h11];
  assign T282 = T283 ? 1'h0 : io_rx_val;
  assign T283 = ! io_rx_val;
  assign T284 = T283 ? 1'h0 : T285;
  assign T285 = io_rx_val ? T286 : 1'h0;
  assign T286 = T287;
  assign T287 = in[5'h10:5'h10];
  assign T288 = T289 ? 1'h0 : io_rx_val;
  assign T289 = ! io_rx_val;
  assign T290 = T289 ? 1'h0 : T291;
  assign T291 = io_rx_val ? T292 : 1'h0;
  assign T292 = T293;
  assign T293 = in[4'hf:4'hf];
  assign T294 = T295 ? 1'h0 : io_rx_val;
  assign T295 = ! io_rx_val;
  assign T296 = T295 ? 1'h0 : T297;
  assign T297 = io_rx_val ? T298 : 1'h0;
  assign T298 = T299;
  assign T299 = in[4'he:4'he];
  assign T300 = T301 ? 1'h0 : io_rx_val;
  assign T301 = ! io_rx_val;
  assign T302 = T301 ? 1'h0 : T303;
  assign T303 = io_rx_val ? T304 : 1'h0;
  assign T304 = T305;
  assign T305 = in[4'hd:4'hd];
  assign T306 = T307 ? 1'h0 : io_rx_val;
  assign T307 = ! io_rx_val;
  assign T308 = T307 ? 1'h0 : T309;
  assign T309 = io_rx_val ? T310 : 1'h0;
  assign T310 = T311;
  assign T311 = in[4'hc:4'hc];
  assign T312 = T313 ? 1'h0 : io_rx_val;
  assign T313 = ! io_rx_val;
  assign T314 = T313 ? 1'h0 : T315;
  assign T315 = io_rx_val ? T316 : 1'h0;
  assign T316 = T317;
  assign T317 = in[4'hb:4'hb];
  assign T318 = T319 ? 1'h0 : io_rx_val;
  assign T319 = ! io_rx_val;
  assign T320 = T319 ? 1'h0 : T321;
  assign T321 = io_rx_val ? T322 : 1'h0;
  assign T322 = T323;
  assign T323 = in[4'ha:4'ha];
  assign T324 = T325 ? 1'h0 : io_rx_val;
  assign T325 = ! io_rx_val;
  assign T326 = T325 ? 1'h0 : T327;
  assign T327 = io_rx_val ? T328 : 1'h0;
  assign T328 = T329;
  assign T329 = in[4'h9:4'h9];
  assign T330 = T331 ? 1'h0 : io_rx_val;
  assign T331 = ! io_rx_val;
  assign T332 = T331 ? 1'h0 : T333;
  assign T333 = io_rx_val ? T334 : 1'h0;
  assign T334 = T335;
  assign T335 = in[4'h8:4'h8];
  assign T336 = T337 ? 1'h0 : io_rx_val;
  assign T337 = ! io_rx_val;
  assign T338 = T337 ? 1'h0 : T339;
  assign T339 = io_rx_val ? T340 : 1'h0;
  assign T340 = T341;
  assign T341 = in[3'h7:3'h7];
  assign T342 = T343 ? 1'h0 : io_rx_val;
  assign T343 = ! io_rx_val;
  assign T344 = T343 ? 1'h0 : T345;
  assign T345 = io_rx_val ? T346 : 1'h0;
  assign T346 = T347;
  assign T347 = in[3'h6:3'h6];
  assign T348 = T349 ? 1'h0 : io_rx_val;
  assign T349 = ! io_rx_val;
  assign T350 = T349 ? 1'h0 : T351;
  assign T351 = io_rx_val ? T352 : 1'h0;
  assign T352 = T353;
  assign T353 = in[3'h5:3'h5];
  assign T354 = T355 ? 1'h0 : io_rx_val;
  assign T355 = ! io_rx_val;
  assign T356 = T355 ? 1'h0 : T357;
  assign T357 = io_rx_val ? T358 : 1'h0;
  assign T358 = T359;
  assign T359 = in[3'h4:3'h4];
  assign T360 = T361 ? 1'h0 : io_rx_val;
  assign T361 = ! io_rx_val;
  assign T362 = T361 ? 1'h0 : T363;
  assign T363 = io_rx_val ? T364 : 1'h0;
  assign T364 = T365;
  assign T365 = in[2'h3:2'h3];
  assign T366 = T367 ? 1'h0 : io_rx_val;
  assign T367 = ! io_rx_val;
  assign T368 = T367 ? 1'h0 : T369;
  assign T369 = io_rx_val ? T370 : 1'h0;
  assign T370 = T371;
  assign T371 = in[2'h2:2'h2];
  assign T372 = T373 ? 1'h0 : io_rx_val;
  assign T373 = ! io_rx_val;
  assign T374 = T373 ? 1'h0 : T375;
  assign T375 = io_rx_val ? T376 : 1'h0;
  assign T376 = T377;
  assign T377 = in[1'h1:1'h1];
  assign T378 = T379 ? 1'h0 : io_rx_val;
  assign T379 = ! io_rx_val;
  assign T380 = T379 ? 1'h0 : T381;
  assign T381 = io_rx_val ? T382 : 1'h0;
  assign T382 = T383;
  assign T383 = in[1'h0:1'h0];
  assign io_tx_val = T384;
  assign T384 = T390 ? 1'h0 : T385;
  assign T385 = R386 == 7'h63;
  assign T387 = T389 ? 7'h0 : T388;
  assign T388 = R386 + 7'h1;
  assign T389 = R386 == 7'h63;
  assign T390 = ! T385;
  assign io_tx_dat_int = T391;
  assign T391 = T390 ? check_out : T392;
  assign T392 = T385 ? check_out : check_out;
  assign T393 = T385 || T390;
  assign T394 = T390 ? T395 : 64'h0;
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = {T398, out_0};
  assign out_0 = Cell_0_io_out;
  assign T398 = {T399, out_1};
  assign out_1 = Cell_1_io_out;
  assign T399 = {T400, out_2};
  assign out_2 = Cell_2_io_out;
  assign T400 = {T401, out_3};
  assign out_3 = Cell_3_io_out;
  assign T401 = {T402, out_4};
  assign out_4 = Cell_4_io_out;
  assign T402 = {T403, out_5};
  assign out_5 = Cell_5_io_out;
  assign T403 = {T404, out_6};
  assign out_6 = Cell_6_io_out;
  assign T404 = {T405, out_7};
  assign out_7 = Cell_7_io_out;
  assign T405 = {T406, out_8};
  assign out_8 = Cell_8_io_out;
  assign T406 = {T407, out_9};
  assign out_9 = Cell_9_io_out;
  assign T407 = {T408, out_10};
  assign out_10 = Cell_10_io_out;
  assign T408 = {T409, out_11};
  assign out_11 = Cell_11_io_out;
  assign T409 = {T410, out_12};
  assign out_12 = Cell_12_io_out;
  assign T410 = {T411, out_13};
  assign out_13 = Cell_13_io_out;
  assign T411 = {T412, out_14};
  assign out_14 = Cell_14_io_out;
  assign T412 = {T413, out_15};
  assign out_15 = Cell_15_io_out;
  assign T413 = {T414, out_16};
  assign out_16 = Cell_16_io_out;
  assign T414 = {T415, out_17};
  assign out_17 = Cell_17_io_out;
  assign T415 = {T416, out_18};
  assign out_18 = Cell_18_io_out;
  assign T416 = {T417, out_19};
  assign out_19 = Cell_19_io_out;
  assign T417 = {T418, out_20};
  assign out_20 = Cell_20_io_out;
  assign T418 = {T419, out_21};
  assign out_21 = Cell_21_io_out;
  assign T419 = {T420, out_22};
  assign out_22 = Cell_22_io_out;
  assign T420 = {T421, out_23};
  assign out_23 = Cell_23_io_out;
  assign T421 = {T422, out_24};
  assign out_24 = Cell_24_io_out;
  assign T422 = {T423, out_25};
  assign out_25 = Cell_25_io_out;
  assign T423 = {T424, out_26};
  assign out_26 = Cell_26_io_out;
  assign T424 = {T425, out_27};
  assign out_27 = Cell_27_io_out;
  assign T425 = {T426, out_28};
  assign out_28 = Cell_28_io_out;
  assign T426 = {T427, out_29};
  assign out_29 = Cell_29_io_out;
  assign T427 = {T428, out_30};
  assign out_30 = Cell_30_io_out;
  assign T428 = {T429, out_31};
  assign out_31 = Cell_31_io_out;
  assign T429 = {T430, out_32};
  assign out_32 = Cell_32_io_out;
  assign T430 = {T431, out_33};
  assign out_33 = Cell_33_io_out;
  assign T431 = {T432, out_34};
  assign out_34 = Cell_34_io_out;
  assign T432 = {T433, out_35};
  assign out_35 = Cell_35_io_out;
  assign T433 = {T434, out_36};
  assign out_36 = Cell_36_io_out;
  assign T434 = {T435, out_37};
  assign out_37 = Cell_37_io_out;
  assign T435 = {T436, out_38};
  assign out_38 = Cell_38_io_out;
  assign T436 = {T437, out_39};
  assign out_39 = Cell_39_io_out;
  assign T437 = {T438, out_40};
  assign out_40 = Cell_40_io_out;
  assign T438 = {T439, out_41};
  assign out_41 = Cell_41_io_out;
  assign T439 = {T440, out_42};
  assign out_42 = Cell_42_io_out;
  assign T440 = {T441, out_43};
  assign out_43 = Cell_43_io_out;
  assign T441 = {T442, out_44};
  assign out_44 = Cell_44_io_out;
  assign T442 = {T443, out_45};
  assign out_45 = Cell_45_io_out;
  assign T443 = {T444, out_46};
  assign out_46 = Cell_46_io_out;
  assign T444 = {T445, out_47};
  assign out_47 = Cell_47_io_out;
  assign T445 = {T446, out_48};
  assign out_48 = Cell_48_io_out;
  assign T446 = {T447, out_49};
  assign out_49 = Cell_49_io_out;
  assign T447 = {T448, out_50};
  assign out_50 = Cell_50_io_out;
  assign T448 = {T449, out_51};
  assign out_51 = Cell_51_io_out;
  assign T449 = {T450, out_52};
  assign out_52 = Cell_52_io_out;
  assign T450 = {T451, out_53};
  assign out_53 = Cell_53_io_out;
  assign T451 = {T452, out_54};
  assign out_54 = Cell_54_io_out;
  assign T452 = {T453, out_55};
  assign out_55 = Cell_55_io_out;
  assign T453 = {T454, out_56};
  assign out_56 = Cell_56_io_out;
  assign T454 = {T455, out_57};
  assign out_57 = Cell_57_io_out;
  assign T455 = {T456, out_58};
  assign out_58 = Cell_58_io_out;
  assign T456 = {T457, out_59};
  assign out_59 = Cell_59_io_out;
  assign T457 = {T458, out_60};
  assign out_60 = Cell_60_io_out;
  assign T458 = {T459, out_61};
  assign out_61 = Cell_61_io_out;
  assign T459 = {out_63, out_62};
  assign out_62 = Cell_62_io_out;
  assign out_63 = Cell_63_io_out;
  assign io_rx_rdy = T460;
  assign T460 = ! is_full;
  assign T461 = T462 || T385;
  assign T462 = T463 || io_rx_val;
  assign T463 = T464 || io_rx_val;
  assign T464 = T465 || io_rx_val;
  assign T465 = T466 || io_rx_val;
  assign T466 = T467 || io_rx_val;
  assign T467 = T468 || io_rx_val;
  assign T468 = T469 || io_rx_val;
  assign T469 = T470 || io_rx_val;
  assign T470 = T471 || io_rx_val;
  assign T471 = T472 || io_rx_val;
  assign T472 = T473 || io_rx_val;
  assign T473 = T474 || io_rx_val;
  assign T474 = T475 || io_rx_val;
  assign T475 = T476 || io_rx_val;
  assign T476 = T477 || io_rx_val;
  assign T477 = T478 || io_rx_val;
  assign T478 = T479 || io_rx_val;
  assign T479 = T480 || io_rx_val;
  assign T480 = T481 || io_rx_val;
  assign T481 = T482 || io_rx_val;
  assign T482 = T483 || io_rx_val;
  assign T483 = T484 || io_rx_val;
  assign T484 = T485 || io_rx_val;
  assign T485 = T486 || io_rx_val;
  assign T486 = T487 || io_rx_val;
  assign T487 = T488 || io_rx_val;
  assign T488 = T489 || io_rx_val;
  assign T489 = T490 || io_rx_val;
  assign T490 = T491 || io_rx_val;
  assign T491 = T492 || io_rx_val;
  assign T492 = T493 || io_rx_val;
  assign T493 = T494 || io_rx_val;
  assign T494 = T495 || io_rx_val;
  assign T495 = T496 || io_rx_val;
  assign T496 = T497 || io_rx_val;
  assign T497 = T498 || io_rx_val;
  assign T498 = T499 || io_rx_val;
  assign T499 = T500 || io_rx_val;
  assign T500 = T501 || io_rx_val;
  assign T501 = T502 || io_rx_val;
  assign T502 = T503 || io_rx_val;
  assign T503 = T504 || io_rx_val;
  assign T504 = T505 || io_rx_val;
  assign T505 = T506 || io_rx_val;
  assign T506 = T507 || io_rx_val;
  assign T507 = T508 || io_rx_val;
  assign T508 = T509 || io_rx_val;
  assign T509 = T510 || io_rx_val;
  assign T510 = T511 || io_rx_val;
  assign T511 = T512 || io_rx_val;
  assign T512 = T513 || io_rx_val;
  assign T513 = T514 || io_rx_val;
  assign T514 = T515 || io_rx_val;
  assign T515 = T516 || io_rx_val;
  assign T516 = T517 || io_rx_val;
  assign T517 = T518 || io_rx_val;
  assign T518 = T519 || io_rx_val;
  assign T519 = T520 || io_rx_val;
  assign T520 = T521 || io_rx_val;
  assign T521 = T522 || io_rx_val;
  assign T522 = T523 || io_rx_val;
  assign T523 = T524 || io_rx_val;
  assign T524 = io_rx_val || io_rx_val;
  assign T525 = T385 ? 1'h0 : 1'h1;
  Cell Cell_0(.clk(clk),
       .io_in( T380 ),
       .io_in_val( T378 ),
       .io_nbrs_0( Cell_63_io_out ),
       .io_nbrs_1( Cell_56_io_out ),
       .io_nbrs_2( Cell_57_io_out ),
       .io_nbrs_3( Cell_7_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_1_io_out ),
       .io_nbrs_6( Cell_15_io_out ),
       .io_nbrs_7( Cell_8_io_out ),
       .io_nbrs_8( Cell_9_io_out ),
       .io_out( Cell_0_io_out )
  );
  Cell Cell_1(.clk(clk),
       .io_in( T374 ),
       .io_in_val( T372 ),
       .io_nbrs_0( Cell_7_io_out ),
       .io_nbrs_1( Cell_0_io_out ),
       .io_nbrs_2( Cell_1_io_out ),
       .io_nbrs_3( Cell_15_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_9_io_out ),
       .io_nbrs_6( Cell_23_io_out ),
       .io_nbrs_7( Cell_16_io_out ),
       .io_nbrs_8( Cell_17_io_out ),
       .io_out( Cell_1_io_out )
  );
  Cell Cell_2(.clk(clk),
       .io_in( T368 ),
       .io_in_val( T366 ),
       .io_nbrs_0( Cell_15_io_out ),
       .io_nbrs_1( Cell_8_io_out ),
       .io_nbrs_2( Cell_9_io_out ),
       .io_nbrs_3( Cell_23_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_17_io_out ),
       .io_nbrs_6( Cell_31_io_out ),
       .io_nbrs_7( Cell_24_io_out ),
       .io_nbrs_8( Cell_25_io_out ),
       .io_out( Cell_2_io_out )
  );
  Cell Cell_3(.clk(clk),
       .io_in( T362 ),
       .io_in_val( T360 ),
       .io_nbrs_0( Cell_23_io_out ),
       .io_nbrs_1( Cell_16_io_out ),
       .io_nbrs_2( Cell_17_io_out ),
       .io_nbrs_3( Cell_31_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_25_io_out ),
       .io_nbrs_6( Cell_39_io_out ),
       .io_nbrs_7( Cell_32_io_out ),
       .io_nbrs_8( Cell_33_io_out ),
       .io_out( Cell_3_io_out )
  );
  Cell Cell_4(.clk(clk),
       .io_in( T356 ),
       .io_in_val( T354 ),
       .io_nbrs_0( Cell_31_io_out ),
       .io_nbrs_1( Cell_24_io_out ),
       .io_nbrs_2( Cell_25_io_out ),
       .io_nbrs_3( Cell_39_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_33_io_out ),
       .io_nbrs_6( Cell_47_io_out ),
       .io_nbrs_7( Cell_40_io_out ),
       .io_nbrs_8( Cell_41_io_out ),
       .io_out( Cell_4_io_out )
  );
  Cell Cell_5(.clk(clk),
       .io_in( T350 ),
       .io_in_val( T348 ),
       .io_nbrs_0( Cell_39_io_out ),
       .io_nbrs_1( Cell_32_io_out ),
       .io_nbrs_2( Cell_33_io_out ),
       .io_nbrs_3( Cell_47_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_41_io_out ),
       .io_nbrs_6( Cell_55_io_out ),
       .io_nbrs_7( Cell_48_io_out ),
       .io_nbrs_8( Cell_49_io_out ),
       .io_out( Cell_5_io_out )
  );
  Cell Cell_6(.clk(clk),
       .io_in( T344 ),
       .io_in_val( T342 ),
       .io_nbrs_0( Cell_47_io_out ),
       .io_nbrs_1( Cell_40_io_out ),
       .io_nbrs_2( Cell_41_io_out ),
       .io_nbrs_3( Cell_55_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_49_io_out ),
       .io_nbrs_6( Cell_63_io_out ),
       .io_nbrs_7( Cell_56_io_out ),
       .io_nbrs_8( Cell_57_io_out ),
       .io_out( Cell_6_io_out )
  );
  Cell Cell_7(.clk(clk),
       .io_in( T338 ),
       .io_in_val( T336 ),
       .io_nbrs_0( Cell_55_io_out ),
       .io_nbrs_1( Cell_48_io_out ),
       .io_nbrs_2( Cell_49_io_out ),
       .io_nbrs_3( Cell_63_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_57_io_out ),
       .io_nbrs_6( Cell_7_io_out ),
       .io_nbrs_7( Cell_0_io_out ),
       .io_nbrs_8( Cell_1_io_out ),
       .io_out( Cell_7_io_out )
  );
  Cell Cell_8(.clk(clk),
       .io_in( T332 ),
       .io_in_val( T330 ),
       .io_nbrs_0( Cell_56_io_out ),
       .io_nbrs_1( Cell_57_io_out ),
       .io_nbrs_2( Cell_58_io_out ),
       .io_nbrs_3( Cell_0_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_2_io_out ),
       .io_nbrs_6( Cell_8_io_out ),
       .io_nbrs_7( Cell_9_io_out ),
       .io_nbrs_8( Cell_10_io_out ),
       .io_out( Cell_8_io_out )
  );
  Cell Cell_9(.clk(clk),
       .io_in( T326 ),
       .io_in_val( T324 ),
       .io_nbrs_0( Cell_0_io_out ),
       .io_nbrs_1( Cell_1_io_out ),
       .io_nbrs_2( Cell_2_io_out ),
       .io_nbrs_3( Cell_8_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_10_io_out ),
       .io_nbrs_6( Cell_16_io_out ),
       .io_nbrs_7( Cell_17_io_out ),
       .io_nbrs_8( Cell_18_io_out ),
       .io_out( Cell_9_io_out )
  );
  Cell Cell_10(.clk(clk),
       .io_in( T320 ),
       .io_in_val( T318 ),
       .io_nbrs_0( Cell_8_io_out ),
       .io_nbrs_1( Cell_9_io_out ),
       .io_nbrs_2( Cell_10_io_out ),
       .io_nbrs_3( Cell_16_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_18_io_out ),
       .io_nbrs_6( Cell_24_io_out ),
       .io_nbrs_7( Cell_25_io_out ),
       .io_nbrs_8( Cell_26_io_out ),
       .io_out( Cell_10_io_out )
  );
  Cell Cell_11(.clk(clk),
       .io_in( T314 ),
       .io_in_val( T312 ),
       .io_nbrs_0( Cell_16_io_out ),
       .io_nbrs_1( Cell_17_io_out ),
       .io_nbrs_2( Cell_18_io_out ),
       .io_nbrs_3( Cell_24_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_26_io_out ),
       .io_nbrs_6( Cell_32_io_out ),
       .io_nbrs_7( Cell_33_io_out ),
       .io_nbrs_8( Cell_34_io_out ),
       .io_out( Cell_11_io_out )
  );
  Cell Cell_12(.clk(clk),
       .io_in( T308 ),
       .io_in_val( T306 ),
       .io_nbrs_0( Cell_24_io_out ),
       .io_nbrs_1( Cell_25_io_out ),
       .io_nbrs_2( Cell_26_io_out ),
       .io_nbrs_3( Cell_32_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_34_io_out ),
       .io_nbrs_6( Cell_40_io_out ),
       .io_nbrs_7( Cell_41_io_out ),
       .io_nbrs_8( Cell_42_io_out ),
       .io_out( Cell_12_io_out )
  );
  Cell Cell_13(.clk(clk),
       .io_in( T302 ),
       .io_in_val( T300 ),
       .io_nbrs_0( Cell_32_io_out ),
       .io_nbrs_1( Cell_33_io_out ),
       .io_nbrs_2( Cell_34_io_out ),
       .io_nbrs_3( Cell_40_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_42_io_out ),
       .io_nbrs_6( Cell_48_io_out ),
       .io_nbrs_7( Cell_49_io_out ),
       .io_nbrs_8( Cell_50_io_out ),
       .io_out( Cell_13_io_out )
  );
  Cell Cell_14(.clk(clk),
       .io_in( T296 ),
       .io_in_val( T294 ),
       .io_nbrs_0( Cell_40_io_out ),
       .io_nbrs_1( Cell_41_io_out ),
       .io_nbrs_2( Cell_42_io_out ),
       .io_nbrs_3( Cell_48_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_50_io_out ),
       .io_nbrs_6( Cell_56_io_out ),
       .io_nbrs_7( Cell_57_io_out ),
       .io_nbrs_8( Cell_58_io_out ),
       .io_out( Cell_14_io_out )
  );
  Cell Cell_15(.clk(clk),
       .io_in( T290 ),
       .io_in_val( T288 ),
       .io_nbrs_0( Cell_48_io_out ),
       .io_nbrs_1( Cell_49_io_out ),
       .io_nbrs_2( Cell_50_io_out ),
       .io_nbrs_3( Cell_56_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_58_io_out ),
       .io_nbrs_6( Cell_0_io_out ),
       .io_nbrs_7( Cell_1_io_out ),
       .io_nbrs_8( Cell_2_io_out ),
       .io_out( Cell_15_io_out )
  );
  Cell Cell_16(.clk(clk),
       .io_in( T284 ),
       .io_in_val( T282 ),
       .io_nbrs_0( Cell_57_io_out ),
       .io_nbrs_1( Cell_58_io_out ),
       .io_nbrs_2( Cell_59_io_out ),
       .io_nbrs_3( Cell_1_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_3_io_out ),
       .io_nbrs_6( Cell_9_io_out ),
       .io_nbrs_7( Cell_10_io_out ),
       .io_nbrs_8( Cell_11_io_out ),
       .io_out( Cell_16_io_out )
  );
  Cell Cell_17(.clk(clk),
       .io_in( T278 ),
       .io_in_val( T276 ),
       .io_nbrs_0( Cell_1_io_out ),
       .io_nbrs_1( Cell_2_io_out ),
       .io_nbrs_2( Cell_3_io_out ),
       .io_nbrs_3( Cell_9_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_11_io_out ),
       .io_nbrs_6( Cell_17_io_out ),
       .io_nbrs_7( Cell_18_io_out ),
       .io_nbrs_8( Cell_19_io_out ),
       .io_out( Cell_17_io_out )
  );
  Cell Cell_18(.clk(clk),
       .io_in( T272 ),
       .io_in_val( T270 ),
       .io_nbrs_0( Cell_9_io_out ),
       .io_nbrs_1( Cell_10_io_out ),
       .io_nbrs_2( Cell_11_io_out ),
       .io_nbrs_3( Cell_17_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_19_io_out ),
       .io_nbrs_6( Cell_25_io_out ),
       .io_nbrs_7( Cell_26_io_out ),
       .io_nbrs_8( Cell_27_io_out ),
       .io_out( Cell_18_io_out )
  );
  Cell Cell_19(.clk(clk),
       .io_in( T266 ),
       .io_in_val( T264 ),
       .io_nbrs_0( Cell_17_io_out ),
       .io_nbrs_1( Cell_18_io_out ),
       .io_nbrs_2( Cell_19_io_out ),
       .io_nbrs_3( Cell_25_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_27_io_out ),
       .io_nbrs_6( Cell_33_io_out ),
       .io_nbrs_7( Cell_34_io_out ),
       .io_nbrs_8( Cell_35_io_out ),
       .io_out( Cell_19_io_out )
  );
  Cell Cell_20(.clk(clk),
       .io_in( T260 ),
       .io_in_val( T258 ),
       .io_nbrs_0( Cell_25_io_out ),
       .io_nbrs_1( Cell_26_io_out ),
       .io_nbrs_2( Cell_27_io_out ),
       .io_nbrs_3( Cell_33_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_35_io_out ),
       .io_nbrs_6( Cell_41_io_out ),
       .io_nbrs_7( Cell_42_io_out ),
       .io_nbrs_8( Cell_43_io_out ),
       .io_out( Cell_20_io_out )
  );
  Cell Cell_21(.clk(clk),
       .io_in( T254 ),
       .io_in_val( T252 ),
       .io_nbrs_0( Cell_33_io_out ),
       .io_nbrs_1( Cell_34_io_out ),
       .io_nbrs_2( Cell_35_io_out ),
       .io_nbrs_3( Cell_41_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_43_io_out ),
       .io_nbrs_6( Cell_49_io_out ),
       .io_nbrs_7( Cell_50_io_out ),
       .io_nbrs_8( Cell_51_io_out ),
       .io_out( Cell_21_io_out )
  );
  Cell Cell_22(.clk(clk),
       .io_in( T248 ),
       .io_in_val( T246 ),
       .io_nbrs_0( Cell_41_io_out ),
       .io_nbrs_1( Cell_42_io_out ),
       .io_nbrs_2( Cell_43_io_out ),
       .io_nbrs_3( Cell_49_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_51_io_out ),
       .io_nbrs_6( Cell_57_io_out ),
       .io_nbrs_7( Cell_58_io_out ),
       .io_nbrs_8( Cell_59_io_out ),
       .io_out( Cell_22_io_out )
  );
  Cell Cell_23(.clk(clk),
       .io_in( T242 ),
       .io_in_val( T240 ),
       .io_nbrs_0( Cell_49_io_out ),
       .io_nbrs_1( Cell_50_io_out ),
       .io_nbrs_2( Cell_51_io_out ),
       .io_nbrs_3( Cell_57_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_59_io_out ),
       .io_nbrs_6( Cell_1_io_out ),
       .io_nbrs_7( Cell_2_io_out ),
       .io_nbrs_8( Cell_3_io_out ),
       .io_out( Cell_23_io_out )
  );
  Cell Cell_24(.clk(clk),
       .io_in( T236 ),
       .io_in_val( T234 ),
       .io_nbrs_0( Cell_58_io_out ),
       .io_nbrs_1( Cell_59_io_out ),
       .io_nbrs_2( Cell_60_io_out ),
       .io_nbrs_3( Cell_2_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_4_io_out ),
       .io_nbrs_6( Cell_10_io_out ),
       .io_nbrs_7( Cell_11_io_out ),
       .io_nbrs_8( Cell_12_io_out ),
       .io_out( Cell_24_io_out )
  );
  Cell Cell_25(.clk(clk),
       .io_in( T230 ),
       .io_in_val( T228 ),
       .io_nbrs_0( Cell_2_io_out ),
       .io_nbrs_1( Cell_3_io_out ),
       .io_nbrs_2( Cell_4_io_out ),
       .io_nbrs_3( Cell_10_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_12_io_out ),
       .io_nbrs_6( Cell_18_io_out ),
       .io_nbrs_7( Cell_19_io_out ),
       .io_nbrs_8( Cell_20_io_out ),
       .io_out( Cell_25_io_out )
  );
  Cell Cell_26(.clk(clk),
       .io_in( T224 ),
       .io_in_val( T222 ),
       .io_nbrs_0( Cell_10_io_out ),
       .io_nbrs_1( Cell_11_io_out ),
       .io_nbrs_2( Cell_12_io_out ),
       .io_nbrs_3( Cell_18_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_20_io_out ),
       .io_nbrs_6( Cell_26_io_out ),
       .io_nbrs_7( Cell_27_io_out ),
       .io_nbrs_8( Cell_28_io_out ),
       .io_out( Cell_26_io_out )
  );
  Cell Cell_27(.clk(clk),
       .io_in( T218 ),
       .io_in_val( T216 ),
       .io_nbrs_0( Cell_18_io_out ),
       .io_nbrs_1( Cell_19_io_out ),
       .io_nbrs_2( Cell_20_io_out ),
       .io_nbrs_3( Cell_26_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_28_io_out ),
       .io_nbrs_6( Cell_34_io_out ),
       .io_nbrs_7( Cell_35_io_out ),
       .io_nbrs_8( Cell_36_io_out ),
       .io_out( Cell_27_io_out )
  );
  Cell Cell_28(.clk(clk),
       .io_in( T212 ),
       .io_in_val( T210 ),
       .io_nbrs_0( Cell_26_io_out ),
       .io_nbrs_1( Cell_27_io_out ),
       .io_nbrs_2( Cell_28_io_out ),
       .io_nbrs_3( Cell_34_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_36_io_out ),
       .io_nbrs_6( Cell_42_io_out ),
       .io_nbrs_7( Cell_43_io_out ),
       .io_nbrs_8( Cell_44_io_out ),
       .io_out( Cell_28_io_out )
  );
  Cell Cell_29(.clk(clk),
       .io_in( T206 ),
       .io_in_val( T204 ),
       .io_nbrs_0( Cell_34_io_out ),
       .io_nbrs_1( Cell_35_io_out ),
       .io_nbrs_2( Cell_36_io_out ),
       .io_nbrs_3( Cell_42_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_44_io_out ),
       .io_nbrs_6( Cell_50_io_out ),
       .io_nbrs_7( Cell_51_io_out ),
       .io_nbrs_8( Cell_52_io_out ),
       .io_out( Cell_29_io_out )
  );
  Cell Cell_30(.clk(clk),
       .io_in( T200 ),
       .io_in_val( T198 ),
       .io_nbrs_0( Cell_42_io_out ),
       .io_nbrs_1( Cell_43_io_out ),
       .io_nbrs_2( Cell_44_io_out ),
       .io_nbrs_3( Cell_50_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_52_io_out ),
       .io_nbrs_6( Cell_58_io_out ),
       .io_nbrs_7( Cell_59_io_out ),
       .io_nbrs_8( Cell_60_io_out ),
       .io_out( Cell_30_io_out )
  );
  Cell Cell_31(.clk(clk),
       .io_in( T194 ),
       .io_in_val( T192 ),
       .io_nbrs_0( Cell_50_io_out ),
       .io_nbrs_1( Cell_51_io_out ),
       .io_nbrs_2( Cell_52_io_out ),
       .io_nbrs_3( Cell_58_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_60_io_out ),
       .io_nbrs_6( Cell_2_io_out ),
       .io_nbrs_7( Cell_3_io_out ),
       .io_nbrs_8( Cell_4_io_out ),
       .io_out( Cell_31_io_out )
  );
  Cell Cell_32(.clk(clk),
       .io_in( T188 ),
       .io_in_val( T186 ),
       .io_nbrs_0( Cell_59_io_out ),
       .io_nbrs_1( Cell_60_io_out ),
       .io_nbrs_2( Cell_61_io_out ),
       .io_nbrs_3( Cell_3_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_5_io_out ),
       .io_nbrs_6( Cell_11_io_out ),
       .io_nbrs_7( Cell_12_io_out ),
       .io_nbrs_8( Cell_13_io_out ),
       .io_out( Cell_32_io_out )
  );
  Cell Cell_33(.clk(clk),
       .io_in( T182 ),
       .io_in_val( T180 ),
       .io_nbrs_0( Cell_3_io_out ),
       .io_nbrs_1( Cell_4_io_out ),
       .io_nbrs_2( Cell_5_io_out ),
       .io_nbrs_3( Cell_11_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_13_io_out ),
       .io_nbrs_6( Cell_19_io_out ),
       .io_nbrs_7( Cell_20_io_out ),
       .io_nbrs_8( Cell_21_io_out ),
       .io_out( Cell_33_io_out )
  );
  Cell Cell_34(.clk(clk),
       .io_in( T176 ),
       .io_in_val( T174 ),
       .io_nbrs_0( Cell_11_io_out ),
       .io_nbrs_1( Cell_12_io_out ),
       .io_nbrs_2( Cell_13_io_out ),
       .io_nbrs_3( Cell_19_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_21_io_out ),
       .io_nbrs_6( Cell_27_io_out ),
       .io_nbrs_7( Cell_28_io_out ),
       .io_nbrs_8( Cell_29_io_out ),
       .io_out( Cell_34_io_out )
  );
  Cell Cell_35(.clk(clk),
       .io_in( T170 ),
       .io_in_val( T168 ),
       .io_nbrs_0( Cell_19_io_out ),
       .io_nbrs_1( Cell_20_io_out ),
       .io_nbrs_2( Cell_21_io_out ),
       .io_nbrs_3( Cell_27_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_29_io_out ),
       .io_nbrs_6( Cell_35_io_out ),
       .io_nbrs_7( Cell_36_io_out ),
       .io_nbrs_8( Cell_37_io_out ),
       .io_out( Cell_35_io_out )
  );
  Cell Cell_36(.clk(clk),
       .io_in( T164 ),
       .io_in_val( T162 ),
       .io_nbrs_0( Cell_27_io_out ),
       .io_nbrs_1( Cell_28_io_out ),
       .io_nbrs_2( Cell_29_io_out ),
       .io_nbrs_3( Cell_35_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_37_io_out ),
       .io_nbrs_6( Cell_43_io_out ),
       .io_nbrs_7( Cell_44_io_out ),
       .io_nbrs_8( Cell_45_io_out ),
       .io_out( Cell_36_io_out )
  );
  Cell Cell_37(.clk(clk),
       .io_in( T158 ),
       .io_in_val( T156 ),
       .io_nbrs_0( Cell_35_io_out ),
       .io_nbrs_1( Cell_36_io_out ),
       .io_nbrs_2( Cell_37_io_out ),
       .io_nbrs_3( Cell_43_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_45_io_out ),
       .io_nbrs_6( Cell_51_io_out ),
       .io_nbrs_7( Cell_52_io_out ),
       .io_nbrs_8( Cell_53_io_out ),
       .io_out( Cell_37_io_out )
  );
  Cell Cell_38(.clk(clk),
       .io_in( T152 ),
       .io_in_val( T150 ),
       .io_nbrs_0( Cell_43_io_out ),
       .io_nbrs_1( Cell_44_io_out ),
       .io_nbrs_2( Cell_45_io_out ),
       .io_nbrs_3( Cell_51_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_53_io_out ),
       .io_nbrs_6( Cell_59_io_out ),
       .io_nbrs_7( Cell_60_io_out ),
       .io_nbrs_8( Cell_61_io_out ),
       .io_out( Cell_38_io_out )
  );
  Cell Cell_39(.clk(clk),
       .io_in( T146 ),
       .io_in_val( T144 ),
       .io_nbrs_0( Cell_51_io_out ),
       .io_nbrs_1( Cell_52_io_out ),
       .io_nbrs_2( Cell_53_io_out ),
       .io_nbrs_3( Cell_59_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_61_io_out ),
       .io_nbrs_6( Cell_3_io_out ),
       .io_nbrs_7( Cell_4_io_out ),
       .io_nbrs_8( Cell_5_io_out ),
       .io_out( Cell_39_io_out )
  );
  Cell Cell_40(.clk(clk),
       .io_in( T140 ),
       .io_in_val( T138 ),
       .io_nbrs_0( Cell_60_io_out ),
       .io_nbrs_1( Cell_61_io_out ),
       .io_nbrs_2( Cell_62_io_out ),
       .io_nbrs_3( Cell_4_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_6_io_out ),
       .io_nbrs_6( Cell_12_io_out ),
       .io_nbrs_7( Cell_13_io_out ),
       .io_nbrs_8( Cell_14_io_out ),
       .io_out( Cell_40_io_out )
  );
  Cell Cell_41(.clk(clk),
       .io_in( T134 ),
       .io_in_val( T132 ),
       .io_nbrs_0( Cell_4_io_out ),
       .io_nbrs_1( Cell_5_io_out ),
       .io_nbrs_2( Cell_6_io_out ),
       .io_nbrs_3( Cell_12_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_14_io_out ),
       .io_nbrs_6( Cell_20_io_out ),
       .io_nbrs_7( Cell_21_io_out ),
       .io_nbrs_8( Cell_22_io_out ),
       .io_out( Cell_41_io_out )
  );
  Cell Cell_42(.clk(clk),
       .io_in( T128 ),
       .io_in_val( T126 ),
       .io_nbrs_0( Cell_12_io_out ),
       .io_nbrs_1( Cell_13_io_out ),
       .io_nbrs_2( Cell_14_io_out ),
       .io_nbrs_3( Cell_20_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_22_io_out ),
       .io_nbrs_6( Cell_28_io_out ),
       .io_nbrs_7( Cell_29_io_out ),
       .io_nbrs_8( Cell_30_io_out ),
       .io_out( Cell_42_io_out )
  );
  Cell Cell_43(.clk(clk),
       .io_in( T122 ),
       .io_in_val( T120 ),
       .io_nbrs_0( Cell_20_io_out ),
       .io_nbrs_1( Cell_21_io_out ),
       .io_nbrs_2( Cell_22_io_out ),
       .io_nbrs_3( Cell_28_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_30_io_out ),
       .io_nbrs_6( Cell_36_io_out ),
       .io_nbrs_7( Cell_37_io_out ),
       .io_nbrs_8( Cell_38_io_out ),
       .io_out( Cell_43_io_out )
  );
  Cell Cell_44(.clk(clk),
       .io_in( T116 ),
       .io_in_val( T114 ),
       .io_nbrs_0( Cell_28_io_out ),
       .io_nbrs_1( Cell_29_io_out ),
       .io_nbrs_2( Cell_30_io_out ),
       .io_nbrs_3( Cell_36_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_38_io_out ),
       .io_nbrs_6( Cell_44_io_out ),
       .io_nbrs_7( Cell_45_io_out ),
       .io_nbrs_8( Cell_46_io_out ),
       .io_out( Cell_44_io_out )
  );
  Cell Cell_45(.clk(clk),
       .io_in( T110 ),
       .io_in_val( T108 ),
       .io_nbrs_0( Cell_36_io_out ),
       .io_nbrs_1( Cell_37_io_out ),
       .io_nbrs_2( Cell_38_io_out ),
       .io_nbrs_3( Cell_44_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_46_io_out ),
       .io_nbrs_6( Cell_52_io_out ),
       .io_nbrs_7( Cell_53_io_out ),
       .io_nbrs_8( Cell_54_io_out ),
       .io_out( Cell_45_io_out )
  );
  Cell Cell_46(.clk(clk),
       .io_in( T104 ),
       .io_in_val( T102 ),
       .io_nbrs_0( Cell_44_io_out ),
       .io_nbrs_1( Cell_45_io_out ),
       .io_nbrs_2( Cell_46_io_out ),
       .io_nbrs_3( Cell_52_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_54_io_out ),
       .io_nbrs_6( Cell_60_io_out ),
       .io_nbrs_7( Cell_61_io_out ),
       .io_nbrs_8( Cell_62_io_out ),
       .io_out( Cell_46_io_out )
  );
  Cell Cell_47(.clk(clk),
       .io_in( T98 ),
       .io_in_val( T96 ),
       .io_nbrs_0( Cell_52_io_out ),
       .io_nbrs_1( Cell_53_io_out ),
       .io_nbrs_2( Cell_54_io_out ),
       .io_nbrs_3( Cell_60_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_62_io_out ),
       .io_nbrs_6( Cell_4_io_out ),
       .io_nbrs_7( Cell_5_io_out ),
       .io_nbrs_8( Cell_6_io_out ),
       .io_out( Cell_47_io_out )
  );
  Cell Cell_48(.clk(clk),
       .io_in( T92 ),
       .io_in_val( T90 ),
       .io_nbrs_0( Cell_61_io_out ),
       .io_nbrs_1( Cell_62_io_out ),
       .io_nbrs_2( Cell_63_io_out ),
       .io_nbrs_3( Cell_5_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_7_io_out ),
       .io_nbrs_6( Cell_13_io_out ),
       .io_nbrs_7( Cell_14_io_out ),
       .io_nbrs_8( Cell_15_io_out ),
       .io_out( Cell_48_io_out )
  );
  Cell Cell_49(.clk(clk),
       .io_in( T86 ),
       .io_in_val( T84 ),
       .io_nbrs_0( Cell_5_io_out ),
       .io_nbrs_1( Cell_6_io_out ),
       .io_nbrs_2( Cell_7_io_out ),
       .io_nbrs_3( Cell_13_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_15_io_out ),
       .io_nbrs_6( Cell_21_io_out ),
       .io_nbrs_7( Cell_22_io_out ),
       .io_nbrs_8( Cell_23_io_out ),
       .io_out( Cell_49_io_out )
  );
  Cell Cell_50(.clk(clk),
       .io_in( T80 ),
       .io_in_val( T78 ),
       .io_nbrs_0( Cell_13_io_out ),
       .io_nbrs_1( Cell_14_io_out ),
       .io_nbrs_2( Cell_15_io_out ),
       .io_nbrs_3( Cell_21_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_23_io_out ),
       .io_nbrs_6( Cell_29_io_out ),
       .io_nbrs_7( Cell_30_io_out ),
       .io_nbrs_8( Cell_31_io_out ),
       .io_out( Cell_50_io_out )
  );
  Cell Cell_51(.clk(clk),
       .io_in( T74 ),
       .io_in_val( T72 ),
       .io_nbrs_0( Cell_21_io_out ),
       .io_nbrs_1( Cell_22_io_out ),
       .io_nbrs_2( Cell_23_io_out ),
       .io_nbrs_3( Cell_29_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_31_io_out ),
       .io_nbrs_6( Cell_37_io_out ),
       .io_nbrs_7( Cell_38_io_out ),
       .io_nbrs_8( Cell_39_io_out ),
       .io_out( Cell_51_io_out )
  );
  Cell Cell_52(.clk(clk),
       .io_in( T68 ),
       .io_in_val( T66 ),
       .io_nbrs_0( Cell_29_io_out ),
       .io_nbrs_1( Cell_30_io_out ),
       .io_nbrs_2( Cell_31_io_out ),
       .io_nbrs_3( Cell_37_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_39_io_out ),
       .io_nbrs_6( Cell_45_io_out ),
       .io_nbrs_7( Cell_46_io_out ),
       .io_nbrs_8( Cell_47_io_out ),
       .io_out( Cell_52_io_out )
  );
  Cell Cell_53(.clk(clk),
       .io_in( T62 ),
       .io_in_val( T60 ),
       .io_nbrs_0( Cell_37_io_out ),
       .io_nbrs_1( Cell_38_io_out ),
       .io_nbrs_2( Cell_39_io_out ),
       .io_nbrs_3( Cell_45_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_47_io_out ),
       .io_nbrs_6( Cell_53_io_out ),
       .io_nbrs_7( Cell_54_io_out ),
       .io_nbrs_8( Cell_55_io_out ),
       .io_out( Cell_53_io_out )
  );
  Cell Cell_54(.clk(clk),
       .io_in( T56 ),
       .io_in_val( T54 ),
       .io_nbrs_0( Cell_45_io_out ),
       .io_nbrs_1( Cell_46_io_out ),
       .io_nbrs_2( Cell_47_io_out ),
       .io_nbrs_3( Cell_53_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_55_io_out ),
       .io_nbrs_6( Cell_61_io_out ),
       .io_nbrs_7( Cell_62_io_out ),
       .io_nbrs_8( Cell_63_io_out ),
       .io_out( Cell_54_io_out )
  );
  Cell Cell_55(.clk(clk),
       .io_in( T50 ),
       .io_in_val( T48 ),
       .io_nbrs_0( Cell_53_io_out ),
       .io_nbrs_1( Cell_54_io_out ),
       .io_nbrs_2( Cell_55_io_out ),
       .io_nbrs_3( Cell_61_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_63_io_out ),
       .io_nbrs_6( Cell_5_io_out ),
       .io_nbrs_7( Cell_6_io_out ),
       .io_nbrs_8( Cell_7_io_out ),
       .io_out( Cell_55_io_out )
  );
  Cell Cell_56(.clk(clk),
       .io_in( T44 ),
       .io_in_val( T42 ),
       .io_nbrs_0( Cell_62_io_out ),
       .io_nbrs_1( Cell_63_io_out ),
       .io_nbrs_2( Cell_56_io_out ),
       .io_nbrs_3( Cell_6_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_0_io_out ),
       .io_nbrs_6( Cell_14_io_out ),
       .io_nbrs_7( Cell_15_io_out ),
       .io_nbrs_8( Cell_8_io_out ),
       .io_out( Cell_56_io_out )
  );
  Cell Cell_57(.clk(clk),
       .io_in( T38 ),
       .io_in_val( T36 ),
       .io_nbrs_0( Cell_6_io_out ),
       .io_nbrs_1( Cell_7_io_out ),
       .io_nbrs_2( Cell_0_io_out ),
       .io_nbrs_3( Cell_14_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_8_io_out ),
       .io_nbrs_6( Cell_22_io_out ),
       .io_nbrs_7( Cell_23_io_out ),
       .io_nbrs_8( Cell_16_io_out ),
       .io_out( Cell_57_io_out )
  );
  Cell Cell_58(.clk(clk),
       .io_in( T32 ),
       .io_in_val( T30 ),
       .io_nbrs_0( Cell_14_io_out ),
       .io_nbrs_1( Cell_15_io_out ),
       .io_nbrs_2( Cell_8_io_out ),
       .io_nbrs_3( Cell_22_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_16_io_out ),
       .io_nbrs_6( Cell_30_io_out ),
       .io_nbrs_7( Cell_31_io_out ),
       .io_nbrs_8( Cell_24_io_out ),
       .io_out( Cell_58_io_out )
  );
  Cell Cell_59(.clk(clk),
       .io_in( T26 ),
       .io_in_val( T24 ),
       .io_nbrs_0( Cell_22_io_out ),
       .io_nbrs_1( Cell_23_io_out ),
       .io_nbrs_2( Cell_16_io_out ),
       .io_nbrs_3( Cell_30_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_24_io_out ),
       .io_nbrs_6( Cell_38_io_out ),
       .io_nbrs_7( Cell_39_io_out ),
       .io_nbrs_8( Cell_32_io_out ),
       .io_out( Cell_59_io_out )
  );
  Cell Cell_60(.clk(clk),
       .io_in( T20 ),
       .io_in_val( T18 ),
       .io_nbrs_0( Cell_30_io_out ),
       .io_nbrs_1( Cell_31_io_out ),
       .io_nbrs_2( Cell_24_io_out ),
       .io_nbrs_3( Cell_38_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_32_io_out ),
       .io_nbrs_6( Cell_46_io_out ),
       .io_nbrs_7( Cell_47_io_out ),
       .io_nbrs_8( Cell_40_io_out ),
       .io_out( Cell_60_io_out )
  );
  Cell Cell_61(.clk(clk),
       .io_in( T14 ),
       .io_in_val( T12 ),
       .io_nbrs_0( Cell_38_io_out ),
       .io_nbrs_1( Cell_39_io_out ),
       .io_nbrs_2( Cell_32_io_out ),
       .io_nbrs_3( Cell_46_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_40_io_out ),
       .io_nbrs_6( Cell_54_io_out ),
       .io_nbrs_7( Cell_55_io_out ),
       .io_nbrs_8( Cell_48_io_out ),
       .io_out( Cell_61_io_out )
  );
  Cell Cell_62(.clk(clk),
       .io_in( T8 ),
       .io_in_val( T6 ),
       .io_nbrs_0( Cell_46_io_out ),
       .io_nbrs_1( Cell_47_io_out ),
       .io_nbrs_2( Cell_40_io_out ),
       .io_nbrs_3( Cell_54_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_48_io_out ),
       .io_nbrs_6( Cell_62_io_out ),
       .io_nbrs_7( Cell_63_io_out ),
       .io_nbrs_8( Cell_56_io_out ),
       .io_out( Cell_62_io_out )
  );
  Cell Cell_63(.clk(clk),
       .io_in( T2 ),
       .io_in_val( T0 ),
       .io_nbrs_0( Cell_54_io_out ),
       .io_nbrs_1( Cell_55_io_out ),
       .io_nbrs_2( Cell_48_io_out ),
       .io_nbrs_3( Cell_62_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_56_io_out ),
       .io_nbrs_6( Cell_6_io_out ),
       .io_nbrs_7( Cell_7_io_out ),
       .io_nbrs_8( Cell_0_io_out ),
       .io_out( Cell_63_io_out )
  );

  always @(posedge clk) begin
    R386 <= reset ? 7'h0 : T387;
    if(reset) begin
      check_out <= 64'h1;
    end else if(T393) begin
      check_out <= T394;
    end
    if(reset) begin
      is_full <= 1'h0;
    end else if(T461) begin
      is_full <= T525;
    end
  end
endmodule

module Controller(input clk, input reset,
    input [63:0] io_rx_dat_int,
    input  io_rx_val,
    output[63:0] io_tx_dat_int,
    output io_tx_val
);

  wire T0;
  wire T1;
  wire Fifo_0_io_deq_val;
  wire Mapper_io_rx_rdy;
  wire T2;
  wire[63:0] Fifo_0_io_deq_dat_int;
  wire[63:0] Mapper_io_tx_dat_int;
  wire T3;
  wire Fifo_1_io_deq_val;
  wire T4;
  wire T5;
  wire T6;
  wire Fifo_1_io_enq_rdy;
  wire Mapper_io_tx_val;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire Fifo_0_io_enq_rdy;
  wire T11;
  wire T12;
  reg[0:0] inCounter;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[63:0] T17;
  wire[63:0] Fifo_1_io_deq_dat_int;

  assign T0 = T2 ? 1'h0 : T1;
  assign T1 = Mapper_io_rx_rdy && Fifo_0_io_deq_val;
  assign T2 = ! T1;
  assign T3 = T4 ? 1'h0 : Fifo_1_io_deq_val;
  assign T4 = ! Fifo_1_io_deq_val;
  assign T5 = T7 ? 1'h0 : T6;
  assign T6 = Mapper_io_tx_val && Fifo_1_io_enq_rdy;
  assign T7 = ! T6;
  assign T8 = T2 ? 1'h0 : T1;
  assign T9 = T16 ? 1'h0 : T10;
  assign T10 = T11 && Fifo_0_io_enq_rdy;
  assign T11 = T12 && io_rx_val;
  assign T12 = 1'h0 == inCounter;
  assign T13 = T15 ? 1'h0 : T14;
  assign T14 = inCounter + 1'h1;
  assign T15 = inCounter == 1'h0;
  assign T16 = ! T10;
  assign io_tx_val = Fifo_1_io_deq_val;
  assign io_tx_dat_int = T17;
  assign T17 = Fifo_1_io_deq_val ? Fifo_1_io_deq_dat_int : 64'h0;
  Fifo_1 Fifo_0(.clk(clk), .reset(reset),
       .io_enq_val( T9 ),
       .io_enq_rdy( Fifo_0_io_enq_rdy ),
       .io_deq_val( Fifo_0_io_deq_val ),
       .io_deq_rdy( T8 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_0_io_deq_dat_int )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enq_val( T5 ),
       .io_enq_rdy( Fifo_1_io_enq_rdy ),
       .io_deq_val( Fifo_1_io_deq_val ),
       .io_deq_rdy( T3 ),
       .io_enq_dat_int( Mapper_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_1_io_deq_dat_int )
  );
  Mapper Mapper(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_0_io_deq_dat_int ),
       .io_rx_val( T0 ),
       .io_rx_rdy( Mapper_io_rx_rdy ),
       .io_tx_dat_int( Mapper_io_tx_dat_int ),
       .io_tx_val( Mapper_io_tx_val )
  );

  always @(posedge clk) begin
    if(reset) begin
      inCounter <= 1'h0;
    end else if(T10) begin
      inCounter <= T13;
    end
  end
endmodule

module MrSimSimulation(input clk, input reset,
    input [63:0] io_enq_dat,
    input  io_enq_val,
    output io_enq_rdy,
    output[63:0] io_deq_dat,
    output io_deq_val,
    input  io_deq_rdy
);

  wire decode_io_tx_val;
  wire[63:0] decode_io_tx_dat_int;
  wire T0;
  wire decode_io_rx_rdy;
  wire Fifo_0_io_deq_val;
  wire[63:0] Fifo_0_io_deq_dat;
  wire Controller_io_tx_val;
  wire[63:0] Controller_io_tx_dat_int;
  wire[63:0] encode_io_tx_dat;
  wire encode_io_tx_val;
  wire T1;
  wire Fifo_1_io_deq_val;
  wire[63:0] Fifo_1_io_deq_dat;
  wire Fifo_0_io_enq_rdy;

  assign T0 = Fifo_0_io_deq_val && decode_io_rx_rdy;
  assign T1 = decode_io_rx_rdy && Fifo_0_io_deq_val;
  assign io_deq_val = Fifo_1_io_deq_val;
  assign io_deq_dat = Fifo_1_io_deq_dat;
  assign io_enq_rdy = Fifo_0_io_enq_rdy;
  Fifo_0 Fifo_0(.clk(clk), .reset(reset),
       .io_enq_val( io_enq_val ),
       .io_enq_rdy( Fifo_0_io_enq_rdy ),
       .io_deq_val( Fifo_0_io_deq_val ),
       .io_deq_rdy( T1 ),
       .io_enq_dat( io_enq_dat ),
       .io_deq_dat( Fifo_0_io_deq_dat )
  );
  Fifo_0 Fifo_1(.clk(clk), .reset(reset),
       .io_enq_val( encode_io_tx_val ),
       //.io_enq_rdy(  )
       .io_deq_val( Fifo_1_io_deq_val ),
       .io_deq_rdy( io_deq_rdy ),
       .io_enq_dat( encode_io_tx_dat ),
       .io_deq_dat( Fifo_1_io_deq_dat )
  );
  encode encode(
       .io_rx_dat_int( Controller_io_tx_dat_int ),
       //.io_rx_rdy(  )
       .io_rx_val( Controller_io_tx_val ),
       .io_tx_dat( encode_io_tx_dat ),
       .io_tx_val( encode_io_tx_val )
  );
  decode decode(
       .io_rx_dat( Fifo_0_io_deq_dat ),
       .io_rx_rdy( decode_io_rx_rdy ),
       .io_rx_val( T0 ),
       .io_tx_dat_int( decode_io_tx_dat_int ),
       .io_tx_val( decode_io_tx_val )
  );
  Controller Controller(.clk(clk), .reset(reset),
       .io_rx_dat_int( decode_io_tx_dat_int ),
       .io_rx_val( decode_io_tx_val ),
       .io_tx_dat_int( Controller_io_tx_dat_int ),
       .io_tx_val( Controller_io_tx_val )
  );
endmodule

