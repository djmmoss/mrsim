module Fifo_0(input clk, input reset,
    input  io_enq_val,
    output io_enq_rdy,
    output io_deq_val,
    input  io_deq_rdy,
    input [63:0] io_enq_dat,
    output[63:0] io_deq_dat
);

  wire[63:0] T0;
  wire[63:0] T1;
  reg [63:0] ram [3:0];
  wire[63:0] T2;
  wire[63:0] T3;
  wire do_enq;
  wire T4;
  reg[0:0] is_full;
  wire is_full_next;
  wire T5;
  wire T6;
  wire do_deq;
  wire T7;
  wire is_empty;
  wire T8;
  reg[3:0] deq_ptr;
  wire[3:0] T9;
  wire[3:0] deq_ptr_inc;
  reg[3:0] enq_ptr;
  wire[3:0] T10;
  wire[3:0] enq_ptr_inc;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;

  assign io_deq_dat = T0;
  assign T0 = do_deq ? T1 : 64'h0;
  assign T1 = ram[T17];
  assign T3 = io_enq_dat;
  assign do_enq = T4 && io_enq_val;
  assign T4 = ! is_full;
  assign is_full_next = T12 ? 1'h1 : T5;
  assign T5 = T6 ? 1'h0 : is_full;
  assign T6 = do_deq && is_full;
  assign do_deq = io_deq_rdy && T7;
  assign T7 = ! is_empty;
  assign is_empty = T11 && T8;
  assign T8 = enq_ptr == deq_ptr;
  assign T9 = do_deq ? deq_ptr_inc : deq_ptr;
  assign deq_ptr_inc = deq_ptr + 4'h1;
  assign T10 = do_enq ? enq_ptr_inc : enq_ptr;
  assign enq_ptr_inc = enq_ptr + 4'h1;
  assign T11 = ! is_full;
  assign T12 = T14 && T13;
  assign T13 = enq_ptr_inc == deq_ptr;
  assign T14 = do_enq && T15;
  assign T15 = ~ do_deq;
  assign T16 = enq_ptr[1'h1:1'h0];
  assign T17 = deq_ptr[1'h1:1'h0];
  assign io_deq_val = T18;
  assign T18 = ! is_empty;
  assign io_enq_rdy = T19;
  assign T19 = ! is_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[T16] <= T3;
    is_full <= reset ? 1'h0 : is_full_next;
    deq_ptr <= reset ? 4'h0 : T9;
    enq_ptr <= reset ? 4'h0 : T10;
  end
endmodule

module encode(
    input [63:0] io_rx_dat_int,
    output io_rx_rdy,
    input  io_rx_val,
    output[63:0] io_tx_dat,
    output io_tx_val
);


  assign io_tx_val = io_rx_val;
  assign io_tx_dat = io_rx_dat_int;
  assign io_rx_rdy = 1'h1;
endmodule

module decode(
    input [63:0] io_rx_dat,
    output io_rx_rdy,
    input  io_rx_val,
    output[63:0] io_tx_dat_int,
    output io_tx_val
);


  assign io_tx_val = io_rx_val;
  assign io_tx_dat_int = io_rx_dat;
  assign io_rx_rdy = 1'h1;
endmodule

module Fifo_1(input clk, input reset,
    input  io_enq_val,
    output io_enq_rdy,
    output io_deq_val,
    input  io_deq_rdy,
    input [63:0] io_enq_dat_int,
    output[63:0] io_deq_dat_int
);

  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [63:0] ram [3:0];
  wire[63:0] T4;
  wire[63:0] T5;
  wire do_enq;
  wire T6;
  reg[0:0] is_full;
  wire is_full_next;
  wire T7;
  wire T8;
  wire do_deq;
  wire T9;
  wire is_empty;
  wire T10;
  reg[3:0] deq_ptr;
  wire[3:0] T11;
  wire[3:0] deq_ptr_inc;
  reg[3:0] enq_ptr;
  wire[3:0] T12;
  wire[3:0] enq_ptr_inc;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;

  assign io_deq_dat_int = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = do_deq ? T2 : 64'h0;
  assign T2 = T3[6'h3f:1'h0];
  assign T3 = ram[T19];
  assign T5 = io_enq_dat_int;
  assign do_enq = T6 && io_enq_val;
  assign T6 = ! is_full;
  assign is_full_next = T14 ? 1'h1 : T7;
  assign T7 = T8 ? 1'h0 : is_full;
  assign T8 = do_deq && is_full;
  assign do_deq = io_deq_rdy && T9;
  assign T9 = ! is_empty;
  assign is_empty = T13 && T10;
  assign T10 = enq_ptr == deq_ptr;
  assign T11 = do_deq ? deq_ptr_inc : deq_ptr;
  assign deq_ptr_inc = deq_ptr + 4'h1;
  assign T12 = do_enq ? enq_ptr_inc : enq_ptr;
  assign enq_ptr_inc = enq_ptr + 4'h1;
  assign T13 = ! is_full;
  assign T14 = T16 && T15;
  assign T15 = enq_ptr_inc == deq_ptr;
  assign T16 = do_enq && T17;
  assign T17 = ~ do_deq;
  assign T18 = enq_ptr[1'h1:1'h0];
  assign T19 = deq_ptr[1'h1:1'h0];
  assign io_deq_val = T20;
  assign T20 = ! is_empty;
  assign io_enq_rdy = T21;
  assign T21 = ! is_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[T18] <= T5;
    is_full <= reset ? 1'h0 : is_full_next;
    deq_ptr <= reset ? 4'h0 : T11;
    enq_ptr <= reset ? 4'h0 : T12;
  end
endmodule

module Cell_0(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;

  assign io_out = isAlive;
  assign T0 = T32 || T1;
  assign T1 = T31 && T2;
  assign T2 = T22 && T3;
  assign T3 = T21 && T4;
  assign T4 = count == 3'h3;
  assign count = 3'h0 + T5;
  assign T5 = 3'h0 + T6;
  assign T6 = 3'h0 + T7;
  assign T7 = 3'h0 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T19 + T10;
  assign T10 = T17 + T11;
  assign T11 = T15 + T12;
  assign T12 = T13 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_8;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_7;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_6;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_5;
  assign T21 = ! isAlive;
  assign T22 = ! T23;
  assign T23 = T26 || T24;
  assign T24 = isAlive && T25;
  assign T25 = 3'h4 <= count;
  assign T26 = T29 || T27;
  assign T27 = isAlive && T28;
  assign T28 = count < 3'h4;
  assign T29 = isAlive && T30;
  assign T30 = count < 3'h2;
  assign T31 = ! io_in_val;
  assign T32 = T36 || T33;
  assign T33 = T31 && T34;
  assign T34 = T35 && T24;
  assign T35 = ! T26;
  assign T36 = T40 || T37;
  assign T37 = T31 && T38;
  assign T38 = T39 && T27;
  assign T39 = ! T29;
  assign T40 = io_in_val || T41;
  assign T41 = T31 && T29;
  assign T42 = T1 ? 1'h1 : T43;
  assign T43 = T33 ? 1'h0 : T44;
  assign T44 = T37 ? 1'h1 : T45;
  assign T45 = T41 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T42;
    end
  end
endmodule

module Cell_1(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;

  assign io_out = isAlive;
  assign T0 = T34 || T1;
  assign T1 = T33 && T2;
  assign T2 = T24 && T3;
  assign T3 = T23 && T4;
  assign T4 = count == 3'h3;
  assign count = 3'h0 + T5;
  assign T5 = 3'h0 + T6;
  assign T6 = 3'h0 + T7;
  assign T7 = T21 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T19 + T10;
  assign T10 = T17 + T11;
  assign T11 = T15 + T12;
  assign T12 = T13 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_8;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_7;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_6;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_5;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_3;
  assign T23 = ! isAlive;
  assign T24 = ! T25;
  assign T25 = T28 || T26;
  assign T26 = isAlive && T27;
  assign T27 = 3'h4 <= count;
  assign T28 = T31 || T29;
  assign T29 = isAlive && T30;
  assign T30 = count < 3'h4;
  assign T31 = isAlive && T32;
  assign T32 = count < 3'h2;
  assign T33 = ! io_in_val;
  assign T34 = T38 || T35;
  assign T35 = T33 && T36;
  assign T36 = T37 && T26;
  assign T37 = ! T28;
  assign T38 = T42 || T39;
  assign T39 = T33 && T40;
  assign T40 = T41 && T29;
  assign T41 = ! T31;
  assign T42 = io_in_val || T43;
  assign T43 = T33 && T31;
  assign T44 = T1 ? 1'h1 : T45;
  assign T45 = T35 ? 1'h0 : T46;
  assign T46 = T39 ? 1'h1 : T47;
  assign T47 = T43 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T44;
    end
  end
endmodule

module Cell_2(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;

  assign io_out = isAlive;
  assign T0 = T36 || T1;
  assign T1 = T35 && T2;
  assign T2 = T26 && T3;
  assign T3 = T25 && T4;
  assign T4 = count == 3'h3;
  assign count = 3'h0 + T5;
  assign T5 = 3'h0 + T6;
  assign T6 = T23 + T7;
  assign T7 = T21 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T19 + T10;
  assign T10 = T17 + T11;
  assign T11 = T15 + T12;
  assign T12 = T13 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_8;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_7;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_6;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_5;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_3;
  assign T23 = {2'h0, T24};
  assign T24 = io_nbrs_2;
  assign T25 = ! isAlive;
  assign T26 = ! T27;
  assign T27 = T30 || T28;
  assign T28 = isAlive && T29;
  assign T29 = 3'h4 <= count;
  assign T30 = T33 || T31;
  assign T31 = isAlive && T32;
  assign T32 = count < 3'h4;
  assign T33 = isAlive && T34;
  assign T34 = count < 3'h2;
  assign T35 = ! io_in_val;
  assign T36 = T40 || T37;
  assign T37 = T35 && T38;
  assign T38 = T39 && T28;
  assign T39 = ! T30;
  assign T40 = T44 || T41;
  assign T41 = T35 && T42;
  assign T42 = T43 && T31;
  assign T43 = ! T33;
  assign T44 = io_in_val || T45;
  assign T45 = T35 && T33;
  assign T46 = T1 ? 1'h1 : T47;
  assign T47 = T37 ? 1'h0 : T48;
  assign T48 = T41 ? 1'h1 : T49;
  assign T49 = T45 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T46;
    end
  end
endmodule

module Cell_3(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;

  assign io_out = isAlive;
  assign T0 = T38 || T1;
  assign T1 = T37 && T2;
  assign T2 = T28 && T3;
  assign T3 = T27 && T4;
  assign T4 = count == 3'h3;
  assign count = 3'h0 + T5;
  assign T5 = T25 + T6;
  assign T6 = T23 + T7;
  assign T7 = T21 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T19 + T10;
  assign T10 = T17 + T11;
  assign T11 = T15 + T12;
  assign T12 = T13 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_8;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_7;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_6;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_5;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_3;
  assign T23 = {2'h0, T24};
  assign T24 = io_nbrs_2;
  assign T25 = {2'h0, T26};
  assign T26 = io_nbrs_1;
  assign T27 = ! isAlive;
  assign T28 = ! T29;
  assign T29 = T32 || T30;
  assign T30 = isAlive && T31;
  assign T31 = 3'h4 <= count;
  assign T32 = T35 || T33;
  assign T33 = isAlive && T34;
  assign T34 = count < 3'h4;
  assign T35 = isAlive && T36;
  assign T36 = count < 3'h2;
  assign T37 = ! io_in_val;
  assign T38 = T42 || T39;
  assign T39 = T37 && T40;
  assign T40 = T41 && T30;
  assign T41 = ! T32;
  assign T42 = T46 || T43;
  assign T43 = T37 && T44;
  assign T44 = T45 && T33;
  assign T45 = ! T35;
  assign T46 = io_in_val || T47;
  assign T47 = T37 && T35;
  assign T48 = T1 ? 1'h1 : T49;
  assign T49 = T39 ? 1'h0 : T50;
  assign T50 = T43 ? 1'h1 : T51;
  assign T51 = T47 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T48;
    end
  end
endmodule

module Cell_4(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;

  assign io_out = isAlive;
  assign T0 = T40 || T1;
  assign T1 = T39 && T2;
  assign T2 = T30 && T3;
  assign T3 = T29 && T4;
  assign T4 = count == 3'h3;
  assign count = T27 + T5;
  assign T5 = T25 + T6;
  assign T6 = T23 + T7;
  assign T7 = T21 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T19 + T10;
  assign T10 = T17 + T11;
  assign T11 = T15 + T12;
  assign T12 = T13 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_8;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_7;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_6;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_5;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_3;
  assign T23 = {2'h0, T24};
  assign T24 = io_nbrs_2;
  assign T25 = {2'h0, T26};
  assign T26 = io_nbrs_1;
  assign T27 = {2'h0, T28};
  assign T28 = io_nbrs_0;
  assign T29 = ! isAlive;
  assign T30 = ! T31;
  assign T31 = T34 || T32;
  assign T32 = isAlive && T33;
  assign T33 = 3'h4 <= count;
  assign T34 = T37 || T35;
  assign T35 = isAlive && T36;
  assign T36 = count < 3'h4;
  assign T37 = isAlive && T38;
  assign T38 = count < 3'h2;
  assign T39 = ! io_in_val;
  assign T40 = T44 || T41;
  assign T41 = T39 && T42;
  assign T42 = T43 && T32;
  assign T43 = ! T34;
  assign T44 = T48 || T45;
  assign T45 = T39 && T46;
  assign T46 = T47 && T35;
  assign T47 = ! T37;
  assign T48 = io_in_val || T49;
  assign T49 = T39 && T37;
  assign T50 = T1 ? 1'h1 : T51;
  assign T51 = T41 ? 1'h0 : T52;
  assign T52 = T45 ? 1'h1 : T53;
  assign T53 = T49 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T50;
    end
  end
endmodule

module Cell_5(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;

  assign io_out = isAlive;
  assign T0 = T38 || T1;
  assign T1 = T37 && T2;
  assign T2 = T28 && T3;
  assign T3 = T27 && T4;
  assign T4 = count == 3'h3;
  assign count = T25 + T5;
  assign T5 = T23 + T6;
  assign T6 = T21 + T7;
  assign T7 = T19 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T17 + T10;
  assign T10 = T15 + T11;
  assign T11 = T13 + T12;
  assign T12 = 3'h0 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_7;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_6;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_5;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_3;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_2;
  assign T23 = {2'h0, T24};
  assign T24 = io_nbrs_1;
  assign T25 = {2'h0, T26};
  assign T26 = io_nbrs_0;
  assign T27 = ! isAlive;
  assign T28 = ! T29;
  assign T29 = T32 || T30;
  assign T30 = isAlive && T31;
  assign T31 = 3'h4 <= count;
  assign T32 = T35 || T33;
  assign T33 = isAlive && T34;
  assign T34 = count < 3'h4;
  assign T35 = isAlive && T36;
  assign T36 = count < 3'h2;
  assign T37 = ! io_in_val;
  assign T38 = T42 || T39;
  assign T39 = T37 && T40;
  assign T40 = T41 && T30;
  assign T41 = ! T32;
  assign T42 = T46 || T43;
  assign T43 = T37 && T44;
  assign T44 = T45 && T33;
  assign T45 = ! T35;
  assign T46 = io_in_val || T47;
  assign T47 = T37 && T35;
  assign T48 = T1 ? 1'h1 : T49;
  assign T49 = T39 ? 1'h0 : T50;
  assign T50 = T43 ? 1'h1 : T51;
  assign T51 = T47 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T48;
    end
  end
endmodule

module Cell_6(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire[2:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;

  assign io_out = isAlive;
  assign T0 = T36 || T1;
  assign T1 = T35 && T2;
  assign T2 = T26 && T3;
  assign T3 = T25 && T4;
  assign T4 = count == 3'h3;
  assign count = T23 + T5;
  assign T5 = T21 + T6;
  assign T6 = T19 + T7;
  assign T7 = T17 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T15 + T10;
  assign T10 = T13 + T11;
  assign T11 = 3'h0 + T12;
  assign T12 = 3'h0 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_6;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_5;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_3;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_2;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_1;
  assign T23 = {2'h0, T24};
  assign T24 = io_nbrs_0;
  assign T25 = ! isAlive;
  assign T26 = ! T27;
  assign T27 = T30 || T28;
  assign T28 = isAlive && T29;
  assign T29 = 3'h4 <= count;
  assign T30 = T33 || T31;
  assign T31 = isAlive && T32;
  assign T32 = count < 3'h4;
  assign T33 = isAlive && T34;
  assign T34 = count < 3'h2;
  assign T35 = ! io_in_val;
  assign T36 = T40 || T37;
  assign T37 = T35 && T38;
  assign T38 = T39 && T28;
  assign T39 = ! T30;
  assign T40 = T44 || T41;
  assign T41 = T35 && T42;
  assign T42 = T43 && T31;
  assign T43 = ! T33;
  assign T44 = io_in_val || T45;
  assign T45 = T35 && T33;
  assign T46 = T1 ? 1'h1 : T47;
  assign T47 = T37 ? 1'h0 : T48;
  assign T48 = T41 ? 1'h1 : T49;
  assign T49 = T45 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T46;
    end
  end
endmodule

module Cell_7(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;

  assign io_out = isAlive;
  assign T0 = T34 || T1;
  assign T1 = T33 && T2;
  assign T2 = T24 && T3;
  assign T3 = T23 && T4;
  assign T4 = count == 3'h3;
  assign count = T21 + T5;
  assign T5 = T19 + T6;
  assign T6 = T17 + T7;
  assign T7 = T15 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = T13 + T10;
  assign T10 = 3'h0 + T11;
  assign T11 = 3'h0 + T12;
  assign T12 = 3'h0 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_5;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_3;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_2;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_1;
  assign T21 = {2'h0, T22};
  assign T22 = io_nbrs_0;
  assign T23 = ! isAlive;
  assign T24 = ! T25;
  assign T25 = T28 || T26;
  assign T26 = isAlive && T27;
  assign T27 = 3'h4 <= count;
  assign T28 = T31 || T29;
  assign T29 = isAlive && T30;
  assign T30 = count < 3'h4;
  assign T31 = isAlive && T32;
  assign T32 = count < 3'h2;
  assign T33 = ! io_in_val;
  assign T34 = T38 || T35;
  assign T35 = T33 && T36;
  assign T36 = T37 && T26;
  assign T37 = ! T28;
  assign T38 = T42 || T39;
  assign T39 = T33 && T40;
  assign T40 = T41 && T29;
  assign T41 = ! T31;
  assign T42 = io_in_val || T43;
  assign T43 = T33 && T31;
  assign T44 = T1 ? 1'h1 : T45;
  assign T45 = T35 ? 1'h0 : T46;
  assign T46 = T39 ? 1'h1 : T47;
  assign T47 = T43 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T44;
    end
  end
endmodule

module Cell_8(input clk,
    input  io_in,
    input  io_in_val,
    input  io_nbrs_0,
    input  io_nbrs_1,
    input  io_nbrs_2,
    input  io_nbrs_3,
    input  io_nbrs_4,
    input  io_nbrs_5,
    input  io_nbrs_6,
    input  io_nbrs_7,
    input  io_nbrs_8,
    output io_out
);

  reg[0:0] isAlive;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire[2:0] count;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;

  assign io_out = isAlive;
  assign T0 = T32 || T1;
  assign T1 = T31 && T2;
  assign T2 = T22 && T3;
  assign T3 = T21 && T4;
  assign T4 = count == 3'h3;
  assign count = T19 + T5;
  assign T5 = T17 + T6;
  assign T6 = T15 + T7;
  assign T7 = T13 + T8;
  assign T8 = 3'h0 + T9;
  assign T9 = 3'h0 + T10;
  assign T10 = 3'h0 + T11;
  assign T11 = 3'h0 + T12;
  assign T12 = 3'h0 + 3'h0;
  assign T13 = {2'h0, T14};
  assign T14 = io_nbrs_3;
  assign T15 = {2'h0, T16};
  assign T16 = io_nbrs_2;
  assign T17 = {2'h0, T18};
  assign T18 = io_nbrs_1;
  assign T19 = {2'h0, T20};
  assign T20 = io_nbrs_0;
  assign T21 = ! isAlive;
  assign T22 = ! T23;
  assign T23 = T26 || T24;
  assign T24 = isAlive && T25;
  assign T25 = 3'h4 <= count;
  assign T26 = T29 || T27;
  assign T27 = isAlive && T28;
  assign T28 = count < 3'h4;
  assign T29 = isAlive && T30;
  assign T30 = count < 3'h2;
  assign T31 = ! io_in_val;
  assign T32 = T36 || T33;
  assign T33 = T31 && T34;
  assign T34 = T35 && T24;
  assign T35 = ! T26;
  assign T36 = T40 || T37;
  assign T37 = T31 && T38;
  assign T38 = T39 && T27;
  assign T39 = ! T29;
  assign T40 = io_in_val || T41;
  assign T41 = T31 && T29;
  assign T42 = T1 ? 1'h1 : T43;
  assign T43 = T33 ? 1'h0 : T44;
  assign T44 = T37 ? 1'h1 : T45;
  assign T45 = T41 ? 1'h0 : io_in;

  always @(posedge clk) begin
    if(T0) begin
      isAlive <= T42;
    end
  end
endmodule

module Mapper(input clk, input reset,
    input [63:0] io_rx_dat_int,
    input  io_rx_val,
    output io_rx_rdy,
    output[63:0] io_tx_dat_int,
    output io_tx_val
);

  wire Cell_62_io_out;
  wire Cell_56_io_out;
  wire Cell_55_io_out;
  wire Cell_54_io_out;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[63:0] in;
  wire Cell_63_io_out;
  wire Cell_61_io_out;
  wire Cell_53_io_out;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire Cell_60_io_out;
  wire Cell_52_io_out;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire Cell_59_io_out;
  wire Cell_51_io_out;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire Cell_58_io_out;
  wire Cell_50_io_out;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire Cell_57_io_out;
  wire Cell_49_io_out;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire Cell_48_io_out;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire Cell_47_io_out;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire Cell_46_io_out;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire Cell_45_io_out;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire Cell_44_io_out;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire Cell_43_io_out;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire Cell_42_io_out;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire Cell_41_io_out;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire Cell_40_io_out;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire Cell_39_io_out;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire Cell_38_io_out;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire Cell_37_io_out;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire Cell_36_io_out;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire Cell_35_io_out;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire Cell_34_io_out;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire Cell_33_io_out;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire Cell_32_io_out;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire Cell_31_io_out;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire Cell_30_io_out;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire Cell_29_io_out;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire Cell_28_io_out;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire Cell_27_io_out;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire Cell_26_io_out;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire Cell_25_io_out;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire Cell_24_io_out;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire Cell_23_io_out;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire Cell_22_io_out;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire Cell_21_io_out;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire Cell_20_io_out;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire Cell_19_io_out;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire Cell_18_io_out;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire Cell_17_io_out;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire Cell_16_io_out;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire Cell_15_io_out;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire Cell_14_io_out;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire Cell_13_io_out;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire Cell_12_io_out;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire Cell_11_io_out;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire Cell_10_io_out;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire Cell_9_io_out;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire Cell_8_io_out;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire Cell_7_io_out;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire Cell_6_io_out;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire Cell_5_io_out;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire Cell_4_io_out;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire Cell_3_io_out;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire Cell_2_io_out;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire Cell_1_io_out;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire Cell_0_io_out;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  reg[4:0] R387;
  wire[4:0] T388;
  wire[4:0] T389;
  wire T390;
  wire T391;
  reg[63:0] check_out;
  wire T392;
  wire T393;
  wire[63:0] T394;
  wire[63:0] T395;
  wire[63:0] T396;
  wire[63:0] T397;
  wire out_0;
  wire[62:0] T398;
  wire out_1;
  wire[61:0] T399;
  wire out_2;
  wire[60:0] T400;
  wire out_3;
  wire[59:0] T401;
  wire out_4;
  wire[58:0] T402;
  wire out_5;
  wire[57:0] T403;
  wire out_6;
  wire[56:0] T404;
  wire out_7;
  wire[55:0] T405;
  wire out_8;
  wire[54:0] T406;
  wire out_9;
  wire[53:0] T407;
  wire out_10;
  wire[52:0] T408;
  wire out_11;
  wire[51:0] T409;
  wire out_12;
  wire[50:0] T410;
  wire out_13;
  wire[49:0] T411;
  wire out_14;
  wire[48:0] T412;
  wire out_15;
  wire[47:0] T413;
  wire out_16;
  wire[46:0] T414;
  wire out_17;
  wire[45:0] T415;
  wire out_18;
  wire[44:0] T416;
  wire out_19;
  wire[43:0] T417;
  wire out_20;
  wire[42:0] T418;
  wire out_21;
  wire[41:0] T419;
  wire out_22;
  wire[40:0] T420;
  wire out_23;
  wire[39:0] T421;
  wire out_24;
  wire[38:0] T422;
  wire out_25;
  wire[37:0] T423;
  wire out_26;
  wire[36:0] T424;
  wire out_27;
  wire[35:0] T425;
  wire out_28;
  wire[34:0] T426;
  wire out_29;
  wire[33:0] T427;
  wire out_30;
  wire[32:0] T428;
  wire out_31;
  wire[31:0] T429;
  wire out_32;
  wire[30:0] T430;
  wire out_33;
  wire[29:0] T431;
  wire out_34;
  wire[28:0] T432;
  wire out_35;
  wire[27:0] T433;
  wire out_36;
  wire[26:0] T434;
  wire out_37;
  wire[25:0] T435;
  wire out_38;
  wire[24:0] T436;
  wire out_39;
  wire[23:0] T437;
  wire out_40;
  wire[22:0] T438;
  wire out_41;
  wire[21:0] T439;
  wire out_42;
  wire[20:0] T440;
  wire out_43;
  wire[19:0] T441;
  wire out_44;
  wire[18:0] T442;
  wire out_45;
  wire[17:0] T443;
  wire out_46;
  wire[16:0] T444;
  wire out_47;
  wire[15:0] T445;
  wire out_48;
  wire[14:0] T446;
  wire out_49;
  wire[13:0] T447;
  wire out_50;
  wire[12:0] T448;
  wire out_51;
  wire[11:0] T449;
  wire out_52;
  wire[10:0] T450;
  wire out_53;
  wire[9:0] T451;
  wire out_54;
  wire[8:0] T452;
  wire out_55;
  wire[7:0] T453;
  wire out_56;
  wire[6:0] T454;
  wire out_57;
  wire[5:0] T455;
  wire out_58;
  wire[4:0] T456;
  wire out_59;
  wire[3:0] T457;
  wire out_60;
  wire[2:0] T458;
  wire out_61;
  wire[1:0] T459;
  wire out_62;
  wire out_63;
  wire[63:0] T460;
  wire[63:0] T461;
  wire[63:0] T462;
  wire[63:0] T463;
  wire T464;
  reg[0:0] is_full;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;

  assign T0 = T1 ? 1'h0 : io_rx_val;
  assign T1 = ! io_rx_val;
  assign T2 = T1 ? 1'h0 : T3;
  assign T3 = io_rx_val ? T4 : 1'h0;
  assign T4 = T5;
  assign T5 = in[6'h3f:6'h3f];
  assign in = io_rx_dat_int;
  assign T6 = T7 ? 1'h0 : io_rx_val;
  assign T7 = ! io_rx_val;
  assign T8 = T7 ? 1'h0 : T9;
  assign T9 = io_rx_val ? T10 : 1'h0;
  assign T10 = T11;
  assign T11 = in[6'h3e:6'h3e];
  assign T12 = T13 ? 1'h0 : io_rx_val;
  assign T13 = ! io_rx_val;
  assign T14 = T13 ? 1'h0 : T15;
  assign T15 = io_rx_val ? T16 : 1'h0;
  assign T16 = T17;
  assign T17 = in[6'h3d:6'h3d];
  assign T18 = T19 ? 1'h0 : io_rx_val;
  assign T19 = ! io_rx_val;
  assign T20 = T19 ? 1'h0 : T21;
  assign T21 = io_rx_val ? T22 : 1'h0;
  assign T22 = T23;
  assign T23 = in[6'h3c:6'h3c];
  assign T24 = T25 ? 1'h0 : io_rx_val;
  assign T25 = ! io_rx_val;
  assign T26 = T25 ? 1'h0 : T27;
  assign T27 = io_rx_val ? T28 : 1'h0;
  assign T28 = T29;
  assign T29 = in[6'h3b:6'h3b];
  assign T30 = T31 ? 1'h0 : io_rx_val;
  assign T31 = ! io_rx_val;
  assign T32 = T31 ? 1'h0 : T33;
  assign T33 = io_rx_val ? T34 : 1'h0;
  assign T34 = T35;
  assign T35 = in[6'h3a:6'h3a];
  assign T36 = T37 ? 1'h0 : io_rx_val;
  assign T37 = ! io_rx_val;
  assign T38 = T37 ? 1'h0 : T39;
  assign T39 = io_rx_val ? T40 : 1'h0;
  assign T40 = T41;
  assign T41 = in[6'h39:6'h39];
  assign T42 = T43 ? 1'h0 : io_rx_val;
  assign T43 = ! io_rx_val;
  assign T44 = T43 ? 1'h0 : T45;
  assign T45 = io_rx_val ? T46 : 1'h0;
  assign T46 = T47;
  assign T47 = in[6'h38:6'h38];
  assign T48 = T49 ? 1'h0 : io_rx_val;
  assign T49 = ! io_rx_val;
  assign T50 = T49 ? 1'h0 : T51;
  assign T51 = io_rx_val ? T52 : 1'h0;
  assign T52 = T53;
  assign T53 = in[6'h37:6'h37];
  assign T54 = T55 ? 1'h0 : io_rx_val;
  assign T55 = ! io_rx_val;
  assign T56 = T55 ? 1'h0 : T57;
  assign T57 = io_rx_val ? T58 : 1'h0;
  assign T58 = T59;
  assign T59 = in[6'h36:6'h36];
  assign T60 = T61 ? 1'h0 : io_rx_val;
  assign T61 = ! io_rx_val;
  assign T62 = T61 ? 1'h0 : T63;
  assign T63 = io_rx_val ? T64 : 1'h0;
  assign T64 = T65;
  assign T65 = in[6'h35:6'h35];
  assign T66 = T67 ? 1'h0 : io_rx_val;
  assign T67 = ! io_rx_val;
  assign T68 = T67 ? 1'h0 : T69;
  assign T69 = io_rx_val ? T70 : 1'h0;
  assign T70 = T71;
  assign T71 = in[6'h34:6'h34];
  assign T72 = T73 ? 1'h0 : io_rx_val;
  assign T73 = ! io_rx_val;
  assign T74 = T73 ? 1'h0 : T75;
  assign T75 = io_rx_val ? T76 : 1'h0;
  assign T76 = T77;
  assign T77 = in[6'h33:6'h33];
  assign T78 = T79 ? 1'h0 : io_rx_val;
  assign T79 = ! io_rx_val;
  assign T80 = T79 ? 1'h0 : T81;
  assign T81 = io_rx_val ? T82 : 1'h0;
  assign T82 = T83;
  assign T83 = in[6'h32:6'h32];
  assign T84 = T85 ? 1'h0 : io_rx_val;
  assign T85 = ! io_rx_val;
  assign T86 = T85 ? 1'h0 : T87;
  assign T87 = io_rx_val ? T88 : 1'h0;
  assign T88 = T89;
  assign T89 = in[6'h31:6'h31];
  assign T90 = T91 ? 1'h0 : io_rx_val;
  assign T91 = ! io_rx_val;
  assign T92 = T91 ? 1'h0 : T93;
  assign T93 = io_rx_val ? T94 : 1'h0;
  assign T94 = T95;
  assign T95 = in[6'h30:6'h30];
  assign T96 = T97 ? 1'h0 : io_rx_val;
  assign T97 = ! io_rx_val;
  assign T98 = T97 ? 1'h0 : T99;
  assign T99 = io_rx_val ? T100 : 1'h0;
  assign T100 = T101;
  assign T101 = in[6'h2f:6'h2f];
  assign T102 = T103 ? 1'h0 : io_rx_val;
  assign T103 = ! io_rx_val;
  assign T104 = T103 ? 1'h0 : T105;
  assign T105 = io_rx_val ? T106 : 1'h0;
  assign T106 = T107;
  assign T107 = in[6'h2e:6'h2e];
  assign T108 = T109 ? 1'h0 : io_rx_val;
  assign T109 = ! io_rx_val;
  assign T110 = T109 ? 1'h0 : T111;
  assign T111 = io_rx_val ? T112 : 1'h0;
  assign T112 = T113;
  assign T113 = in[6'h2d:6'h2d];
  assign T114 = T115 ? 1'h0 : io_rx_val;
  assign T115 = ! io_rx_val;
  assign T116 = T115 ? 1'h0 : T117;
  assign T117 = io_rx_val ? T118 : 1'h0;
  assign T118 = T119;
  assign T119 = in[6'h2c:6'h2c];
  assign T120 = T121 ? 1'h0 : io_rx_val;
  assign T121 = ! io_rx_val;
  assign T122 = T121 ? 1'h0 : T123;
  assign T123 = io_rx_val ? T124 : 1'h0;
  assign T124 = T125;
  assign T125 = in[6'h2b:6'h2b];
  assign T126 = T127 ? 1'h0 : io_rx_val;
  assign T127 = ! io_rx_val;
  assign T128 = T127 ? 1'h0 : T129;
  assign T129 = io_rx_val ? T130 : 1'h0;
  assign T130 = T131;
  assign T131 = in[6'h2a:6'h2a];
  assign T132 = T133 ? 1'h0 : io_rx_val;
  assign T133 = ! io_rx_val;
  assign T134 = T133 ? 1'h0 : T135;
  assign T135 = io_rx_val ? T136 : 1'h0;
  assign T136 = T137;
  assign T137 = in[6'h29:6'h29];
  assign T138 = T139 ? 1'h0 : io_rx_val;
  assign T139 = ! io_rx_val;
  assign T140 = T139 ? 1'h0 : T141;
  assign T141 = io_rx_val ? T142 : 1'h0;
  assign T142 = T143;
  assign T143 = in[6'h28:6'h28];
  assign T144 = T145 ? 1'h0 : io_rx_val;
  assign T145 = ! io_rx_val;
  assign T146 = T145 ? 1'h0 : T147;
  assign T147 = io_rx_val ? T148 : 1'h0;
  assign T148 = T149;
  assign T149 = in[6'h27:6'h27];
  assign T150 = T151 ? 1'h0 : io_rx_val;
  assign T151 = ! io_rx_val;
  assign T152 = T151 ? 1'h0 : T153;
  assign T153 = io_rx_val ? T154 : 1'h0;
  assign T154 = T155;
  assign T155 = in[6'h26:6'h26];
  assign T156 = T157 ? 1'h0 : io_rx_val;
  assign T157 = ! io_rx_val;
  assign T158 = T157 ? 1'h0 : T159;
  assign T159 = io_rx_val ? T160 : 1'h0;
  assign T160 = T161;
  assign T161 = in[6'h25:6'h25];
  assign T162 = T163 ? 1'h0 : io_rx_val;
  assign T163 = ! io_rx_val;
  assign T164 = T163 ? 1'h0 : T165;
  assign T165 = io_rx_val ? T166 : 1'h0;
  assign T166 = T167;
  assign T167 = in[6'h24:6'h24];
  assign T168 = T169 ? 1'h0 : io_rx_val;
  assign T169 = ! io_rx_val;
  assign T170 = T169 ? 1'h0 : T171;
  assign T171 = io_rx_val ? T172 : 1'h0;
  assign T172 = T173;
  assign T173 = in[6'h23:6'h23];
  assign T174 = T175 ? 1'h0 : io_rx_val;
  assign T175 = ! io_rx_val;
  assign T176 = T175 ? 1'h0 : T177;
  assign T177 = io_rx_val ? T178 : 1'h0;
  assign T178 = T179;
  assign T179 = in[6'h22:6'h22];
  assign T180 = T181 ? 1'h0 : io_rx_val;
  assign T181 = ! io_rx_val;
  assign T182 = T181 ? 1'h0 : T183;
  assign T183 = io_rx_val ? T184 : 1'h0;
  assign T184 = T185;
  assign T185 = in[6'h21:6'h21];
  assign T186 = T187 ? 1'h0 : io_rx_val;
  assign T187 = ! io_rx_val;
  assign T188 = T187 ? 1'h0 : T189;
  assign T189 = io_rx_val ? T190 : 1'h0;
  assign T190 = T191;
  assign T191 = in[6'h20:6'h20];
  assign T192 = T193 ? 1'h0 : io_rx_val;
  assign T193 = ! io_rx_val;
  assign T194 = T193 ? 1'h0 : T195;
  assign T195 = io_rx_val ? T196 : 1'h0;
  assign T196 = T197;
  assign T197 = in[5'h1f:5'h1f];
  assign T198 = T199 ? 1'h0 : io_rx_val;
  assign T199 = ! io_rx_val;
  assign T200 = T199 ? 1'h0 : T201;
  assign T201 = io_rx_val ? T202 : 1'h0;
  assign T202 = T203;
  assign T203 = in[5'h1e:5'h1e];
  assign T204 = T205 ? 1'h0 : io_rx_val;
  assign T205 = ! io_rx_val;
  assign T206 = T205 ? 1'h0 : T207;
  assign T207 = io_rx_val ? T208 : 1'h0;
  assign T208 = T209;
  assign T209 = in[5'h1d:5'h1d];
  assign T210 = T211 ? 1'h0 : io_rx_val;
  assign T211 = ! io_rx_val;
  assign T212 = T211 ? 1'h0 : T213;
  assign T213 = io_rx_val ? T214 : 1'h0;
  assign T214 = T215;
  assign T215 = in[5'h1c:5'h1c];
  assign T216 = T217 ? 1'h0 : io_rx_val;
  assign T217 = ! io_rx_val;
  assign T218 = T217 ? 1'h0 : T219;
  assign T219 = io_rx_val ? T220 : 1'h0;
  assign T220 = T221;
  assign T221 = in[5'h1b:5'h1b];
  assign T222 = T223 ? 1'h0 : io_rx_val;
  assign T223 = ! io_rx_val;
  assign T224 = T223 ? 1'h0 : T225;
  assign T225 = io_rx_val ? T226 : 1'h0;
  assign T226 = T227;
  assign T227 = in[5'h1a:5'h1a];
  assign T228 = T229 ? 1'h0 : io_rx_val;
  assign T229 = ! io_rx_val;
  assign T230 = T229 ? 1'h0 : T231;
  assign T231 = io_rx_val ? T232 : 1'h0;
  assign T232 = T233;
  assign T233 = in[5'h19:5'h19];
  assign T234 = T235 ? 1'h0 : io_rx_val;
  assign T235 = ! io_rx_val;
  assign T236 = T235 ? 1'h0 : T237;
  assign T237 = io_rx_val ? T238 : 1'h0;
  assign T238 = T239;
  assign T239 = in[5'h18:5'h18];
  assign T240 = T241 ? 1'h0 : io_rx_val;
  assign T241 = ! io_rx_val;
  assign T242 = T241 ? 1'h0 : T243;
  assign T243 = io_rx_val ? T244 : 1'h0;
  assign T244 = T245;
  assign T245 = in[5'h17:5'h17];
  assign T246 = T247 ? 1'h0 : io_rx_val;
  assign T247 = ! io_rx_val;
  assign T248 = T247 ? 1'h0 : T249;
  assign T249 = io_rx_val ? T250 : 1'h0;
  assign T250 = T251;
  assign T251 = in[5'h16:5'h16];
  assign T252 = T253 ? 1'h0 : io_rx_val;
  assign T253 = ! io_rx_val;
  assign T254 = T253 ? 1'h0 : T255;
  assign T255 = io_rx_val ? T256 : 1'h0;
  assign T256 = T257;
  assign T257 = in[5'h15:5'h15];
  assign T258 = T259 ? 1'h0 : io_rx_val;
  assign T259 = ! io_rx_val;
  assign T260 = T259 ? 1'h0 : T261;
  assign T261 = io_rx_val ? T262 : 1'h0;
  assign T262 = T263;
  assign T263 = in[5'h14:5'h14];
  assign T264 = T265 ? 1'h0 : io_rx_val;
  assign T265 = ! io_rx_val;
  assign T266 = T265 ? 1'h0 : T267;
  assign T267 = io_rx_val ? T268 : 1'h0;
  assign T268 = T269;
  assign T269 = in[5'h13:5'h13];
  assign T270 = T271 ? 1'h0 : io_rx_val;
  assign T271 = ! io_rx_val;
  assign T272 = T271 ? 1'h0 : T273;
  assign T273 = io_rx_val ? T274 : 1'h0;
  assign T274 = T275;
  assign T275 = in[5'h12:5'h12];
  assign T276 = T277 ? 1'h0 : io_rx_val;
  assign T277 = ! io_rx_val;
  assign T278 = T277 ? 1'h0 : T279;
  assign T279 = io_rx_val ? T280 : 1'h0;
  assign T280 = T281;
  assign T281 = in[5'h11:5'h11];
  assign T282 = T283 ? 1'h0 : io_rx_val;
  assign T283 = ! io_rx_val;
  assign T284 = T283 ? 1'h0 : T285;
  assign T285 = io_rx_val ? T286 : 1'h0;
  assign T286 = T287;
  assign T287 = in[5'h10:5'h10];
  assign T288 = T289 ? 1'h0 : io_rx_val;
  assign T289 = ! io_rx_val;
  assign T290 = T289 ? 1'h0 : T291;
  assign T291 = io_rx_val ? T292 : 1'h0;
  assign T292 = T293;
  assign T293 = in[4'hf:4'hf];
  assign T294 = T295 ? 1'h0 : io_rx_val;
  assign T295 = ! io_rx_val;
  assign T296 = T295 ? 1'h0 : T297;
  assign T297 = io_rx_val ? T298 : 1'h0;
  assign T298 = T299;
  assign T299 = in[4'he:4'he];
  assign T300 = T301 ? 1'h0 : io_rx_val;
  assign T301 = ! io_rx_val;
  assign T302 = T301 ? 1'h0 : T303;
  assign T303 = io_rx_val ? T304 : 1'h0;
  assign T304 = T305;
  assign T305 = in[4'hd:4'hd];
  assign T306 = T307 ? 1'h0 : io_rx_val;
  assign T307 = ! io_rx_val;
  assign T308 = T307 ? 1'h0 : T309;
  assign T309 = io_rx_val ? T310 : 1'h0;
  assign T310 = T311;
  assign T311 = in[4'hc:4'hc];
  assign T312 = T313 ? 1'h0 : io_rx_val;
  assign T313 = ! io_rx_val;
  assign T314 = T313 ? 1'h0 : T315;
  assign T315 = io_rx_val ? T316 : 1'h0;
  assign T316 = T317;
  assign T317 = in[4'hb:4'hb];
  assign T318 = T319 ? 1'h0 : io_rx_val;
  assign T319 = ! io_rx_val;
  assign T320 = T319 ? 1'h0 : T321;
  assign T321 = io_rx_val ? T322 : 1'h0;
  assign T322 = T323;
  assign T323 = in[4'ha:4'ha];
  assign T324 = T325 ? 1'h0 : io_rx_val;
  assign T325 = ! io_rx_val;
  assign T326 = T325 ? 1'h0 : T327;
  assign T327 = io_rx_val ? T328 : 1'h0;
  assign T328 = T329;
  assign T329 = in[4'h9:4'h9];
  assign T330 = T331 ? 1'h0 : io_rx_val;
  assign T331 = ! io_rx_val;
  assign T332 = T331 ? 1'h0 : T333;
  assign T333 = io_rx_val ? T334 : 1'h0;
  assign T334 = T335;
  assign T335 = in[4'h8:4'h8];
  assign T336 = T337 ? 1'h0 : io_rx_val;
  assign T337 = ! io_rx_val;
  assign T338 = T337 ? 1'h0 : T339;
  assign T339 = io_rx_val ? T340 : 1'h0;
  assign T340 = T341;
  assign T341 = in[3'h7:3'h7];
  assign T342 = T343 ? 1'h0 : io_rx_val;
  assign T343 = ! io_rx_val;
  assign T344 = T343 ? 1'h0 : T345;
  assign T345 = io_rx_val ? T346 : 1'h0;
  assign T346 = T347;
  assign T347 = in[3'h6:3'h6];
  assign T348 = T349 ? 1'h0 : io_rx_val;
  assign T349 = ! io_rx_val;
  assign T350 = T349 ? 1'h0 : T351;
  assign T351 = io_rx_val ? T352 : 1'h0;
  assign T352 = T353;
  assign T353 = in[3'h5:3'h5];
  assign T354 = T355 ? 1'h0 : io_rx_val;
  assign T355 = ! io_rx_val;
  assign T356 = T355 ? 1'h0 : T357;
  assign T357 = io_rx_val ? T358 : 1'h0;
  assign T358 = T359;
  assign T359 = in[3'h4:3'h4];
  assign T360 = T361 ? 1'h0 : io_rx_val;
  assign T361 = ! io_rx_val;
  assign T362 = T361 ? 1'h0 : T363;
  assign T363 = io_rx_val ? T364 : 1'h0;
  assign T364 = T365;
  assign T365 = in[2'h3:2'h3];
  assign T366 = T367 ? 1'h0 : io_rx_val;
  assign T367 = ! io_rx_val;
  assign T368 = T367 ? 1'h0 : T369;
  assign T369 = io_rx_val ? T370 : 1'h0;
  assign T370 = T371;
  assign T371 = in[2'h2:2'h2];
  assign T372 = T373 ? 1'h0 : io_rx_val;
  assign T373 = ! io_rx_val;
  assign T374 = T373 ? 1'h0 : T375;
  assign T375 = io_rx_val ? T376 : 1'h0;
  assign T376 = T377;
  assign T377 = in[1'h1:1'h1];
  assign T378 = T379 ? 1'h0 : io_rx_val;
  assign T379 = ! io_rx_val;
  assign T380 = T379 ? 1'h0 : T381;
  assign T381 = io_rx_val ? T382 : 1'h0;
  assign T382 = T383;
  assign T383 = in[1'h0:1'h0];
  assign io_tx_val = T384;
  assign T384 = T393 ? 1'h0 : T385;
  assign T385 = T391 || T386;
  assign T386 = R387 == 5'h13;
  assign T388 = T390 ? 5'h0 : T389;
  assign T389 = R387 + 5'h1;
  assign T390 = R387 == 5'h14;
  assign T391 = T460 == check_out;
  assign T392 = T385 || T393;
  assign T393 = ! T385;
  assign T394 = T393 ? T395 : 64'h0;
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = {T398, out_0};
  assign out_0 = Cell_0_io_out;
  assign T398 = {T399, out_1};
  assign out_1 = Cell_1_io_out;
  assign T399 = {T400, out_2};
  assign out_2 = Cell_2_io_out;
  assign T400 = {T401, out_3};
  assign out_3 = Cell_3_io_out;
  assign T401 = {T402, out_4};
  assign out_4 = Cell_4_io_out;
  assign T402 = {T403, out_5};
  assign out_5 = Cell_5_io_out;
  assign T403 = {T404, out_6};
  assign out_6 = Cell_6_io_out;
  assign T404 = {T405, out_7};
  assign out_7 = Cell_7_io_out;
  assign T405 = {T406, out_8};
  assign out_8 = Cell_8_io_out;
  assign T406 = {T407, out_9};
  assign out_9 = Cell_9_io_out;
  assign T407 = {T408, out_10};
  assign out_10 = Cell_10_io_out;
  assign T408 = {T409, out_11};
  assign out_11 = Cell_11_io_out;
  assign T409 = {T410, out_12};
  assign out_12 = Cell_12_io_out;
  assign T410 = {T411, out_13};
  assign out_13 = Cell_13_io_out;
  assign T411 = {T412, out_14};
  assign out_14 = Cell_14_io_out;
  assign T412 = {T413, out_15};
  assign out_15 = Cell_15_io_out;
  assign T413 = {T414, out_16};
  assign out_16 = Cell_16_io_out;
  assign T414 = {T415, out_17};
  assign out_17 = Cell_17_io_out;
  assign T415 = {T416, out_18};
  assign out_18 = Cell_18_io_out;
  assign T416 = {T417, out_19};
  assign out_19 = Cell_19_io_out;
  assign T417 = {T418, out_20};
  assign out_20 = Cell_20_io_out;
  assign T418 = {T419, out_21};
  assign out_21 = Cell_21_io_out;
  assign T419 = {T420, out_22};
  assign out_22 = Cell_22_io_out;
  assign T420 = {T421, out_23};
  assign out_23 = Cell_23_io_out;
  assign T421 = {T422, out_24};
  assign out_24 = Cell_24_io_out;
  assign T422 = {T423, out_25};
  assign out_25 = Cell_25_io_out;
  assign T423 = {T424, out_26};
  assign out_26 = Cell_26_io_out;
  assign T424 = {T425, out_27};
  assign out_27 = Cell_27_io_out;
  assign T425 = {T426, out_28};
  assign out_28 = Cell_28_io_out;
  assign T426 = {T427, out_29};
  assign out_29 = Cell_29_io_out;
  assign T427 = {T428, out_30};
  assign out_30 = Cell_30_io_out;
  assign T428 = {T429, out_31};
  assign out_31 = Cell_31_io_out;
  assign T429 = {T430, out_32};
  assign out_32 = Cell_32_io_out;
  assign T430 = {T431, out_33};
  assign out_33 = Cell_33_io_out;
  assign T431 = {T432, out_34};
  assign out_34 = Cell_34_io_out;
  assign T432 = {T433, out_35};
  assign out_35 = Cell_35_io_out;
  assign T433 = {T434, out_36};
  assign out_36 = Cell_36_io_out;
  assign T434 = {T435, out_37};
  assign out_37 = Cell_37_io_out;
  assign T435 = {T436, out_38};
  assign out_38 = Cell_38_io_out;
  assign T436 = {T437, out_39};
  assign out_39 = Cell_39_io_out;
  assign T437 = {T438, out_40};
  assign out_40 = Cell_40_io_out;
  assign T438 = {T439, out_41};
  assign out_41 = Cell_41_io_out;
  assign T439 = {T440, out_42};
  assign out_42 = Cell_42_io_out;
  assign T440 = {T441, out_43};
  assign out_43 = Cell_43_io_out;
  assign T441 = {T442, out_44};
  assign out_44 = Cell_44_io_out;
  assign T442 = {T443, out_45};
  assign out_45 = Cell_45_io_out;
  assign T443 = {T444, out_46};
  assign out_46 = Cell_46_io_out;
  assign T444 = {T445, out_47};
  assign out_47 = Cell_47_io_out;
  assign T445 = {T446, out_48};
  assign out_48 = Cell_48_io_out;
  assign T446 = {T447, out_49};
  assign out_49 = Cell_49_io_out;
  assign T447 = {T448, out_50};
  assign out_50 = Cell_50_io_out;
  assign T448 = {T449, out_51};
  assign out_51 = Cell_51_io_out;
  assign T449 = {T450, out_52};
  assign out_52 = Cell_52_io_out;
  assign T450 = {T451, out_53};
  assign out_53 = Cell_53_io_out;
  assign T451 = {T452, out_54};
  assign out_54 = Cell_54_io_out;
  assign T452 = {T453, out_55};
  assign out_55 = Cell_55_io_out;
  assign T453 = {T454, out_56};
  assign out_56 = Cell_56_io_out;
  assign T454 = {T455, out_57};
  assign out_57 = Cell_57_io_out;
  assign T455 = {T456, out_58};
  assign out_58 = Cell_58_io_out;
  assign T456 = {T457, out_59};
  assign out_59 = Cell_59_io_out;
  assign T457 = {T458, out_60};
  assign out_60 = Cell_60_io_out;
  assign T458 = {T459, out_61};
  assign out_61 = Cell_61_io_out;
  assign T459 = {out_63, out_62};
  assign out_62 = Cell_62_io_out;
  assign out_63 = Cell_63_io_out;
  assign T460 = T461;
  assign T461 = T397;
  assign io_tx_dat_int = T462;
  assign T462 = T393 ? check_out : T463;
  assign T463 = T385 ? check_out : check_out;
  assign io_rx_rdy = T464;
  assign T464 = ! is_full;
  assign T465 = T466 || T385;
  assign T466 = T467 || io_rx_val;
  assign T467 = T468 || io_rx_val;
  assign T468 = T469 || io_rx_val;
  assign T469 = T470 || io_rx_val;
  assign T470 = T471 || io_rx_val;
  assign T471 = T472 || io_rx_val;
  assign T472 = T473 || io_rx_val;
  assign T473 = T474 || io_rx_val;
  assign T474 = T475 || io_rx_val;
  assign T475 = T476 || io_rx_val;
  assign T476 = T477 || io_rx_val;
  assign T477 = T478 || io_rx_val;
  assign T478 = T479 || io_rx_val;
  assign T479 = T480 || io_rx_val;
  assign T480 = T481 || io_rx_val;
  assign T481 = T482 || io_rx_val;
  assign T482 = T483 || io_rx_val;
  assign T483 = T484 || io_rx_val;
  assign T484 = T485 || io_rx_val;
  assign T485 = T486 || io_rx_val;
  assign T486 = T487 || io_rx_val;
  assign T487 = T488 || io_rx_val;
  assign T488 = T489 || io_rx_val;
  assign T489 = T490 || io_rx_val;
  assign T490 = T491 || io_rx_val;
  assign T491 = T492 || io_rx_val;
  assign T492 = T493 || io_rx_val;
  assign T493 = T494 || io_rx_val;
  assign T494 = T495 || io_rx_val;
  assign T495 = T496 || io_rx_val;
  assign T496 = T497 || io_rx_val;
  assign T497 = T498 || io_rx_val;
  assign T498 = T499 || io_rx_val;
  assign T499 = T500 || io_rx_val;
  assign T500 = T501 || io_rx_val;
  assign T501 = T502 || io_rx_val;
  assign T502 = T503 || io_rx_val;
  assign T503 = T504 || io_rx_val;
  assign T504 = T505 || io_rx_val;
  assign T505 = T506 || io_rx_val;
  assign T506 = T507 || io_rx_val;
  assign T507 = T508 || io_rx_val;
  assign T508 = T509 || io_rx_val;
  assign T509 = T510 || io_rx_val;
  assign T510 = T511 || io_rx_val;
  assign T511 = T512 || io_rx_val;
  assign T512 = T513 || io_rx_val;
  assign T513 = T514 || io_rx_val;
  assign T514 = T515 || io_rx_val;
  assign T515 = T516 || io_rx_val;
  assign T516 = T517 || io_rx_val;
  assign T517 = T518 || io_rx_val;
  assign T518 = T519 || io_rx_val;
  assign T519 = T520 || io_rx_val;
  assign T520 = T521 || io_rx_val;
  assign T521 = T522 || io_rx_val;
  assign T522 = T523 || io_rx_val;
  assign T523 = T524 || io_rx_val;
  assign T524 = T525 || io_rx_val;
  assign T525 = T526 || io_rx_val;
  assign T526 = T527 || io_rx_val;
  assign T527 = T528 || io_rx_val;
  assign T528 = io_rx_val || io_rx_val;
  assign T529 = T385 ? 1'h0 : 1'h1;
  Cell_0 Cell_0(.clk(clk),
       .io_in( T380 ),
       .io_in_val( T378 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( 1'h0 ),
       .io_nbrs_3( 1'h0 ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_1_io_out ),
       .io_nbrs_6( Cell_7_io_out ),
       .io_nbrs_7( Cell_8_io_out ),
       .io_nbrs_8( Cell_9_io_out ),
       .io_out( Cell_0_io_out )
  );
  Cell_1 Cell_1(.clk(clk),
       .io_in( T374 ),
       .io_in_val( T372 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( 1'h0 ),
       .io_nbrs_3( Cell_0_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_2_io_out ),
       .io_nbrs_6( Cell_8_io_out ),
       .io_nbrs_7( Cell_9_io_out ),
       .io_nbrs_8( Cell_10_io_out ),
       .io_out( Cell_1_io_out )
  );
  Cell_1 Cell_2(.clk(clk),
       .io_in( T368 ),
       .io_in_val( T366 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( 1'h0 ),
       .io_nbrs_3( Cell_1_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_3_io_out ),
       .io_nbrs_6( Cell_9_io_out ),
       .io_nbrs_7( Cell_10_io_out ),
       .io_nbrs_8( Cell_11_io_out ),
       .io_out( Cell_2_io_out )
  );
  Cell_1 Cell_3(.clk(clk),
       .io_in( T362 ),
       .io_in_val( T360 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( 1'h0 ),
       .io_nbrs_3( Cell_2_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_4_io_out ),
       .io_nbrs_6( Cell_10_io_out ),
       .io_nbrs_7( Cell_11_io_out ),
       .io_nbrs_8( Cell_12_io_out ),
       .io_out( Cell_3_io_out )
  );
  Cell_1 Cell_4(.clk(clk),
       .io_in( T356 ),
       .io_in_val( T354 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( 1'h0 ),
       .io_nbrs_3( Cell_3_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_5_io_out ),
       .io_nbrs_6( Cell_11_io_out ),
       .io_nbrs_7( Cell_12_io_out ),
       .io_nbrs_8( Cell_13_io_out ),
       .io_out( Cell_4_io_out )
  );
  Cell_1 Cell_5(.clk(clk),
       .io_in( T350 ),
       .io_in_val( T348 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( 1'h0 ),
       .io_nbrs_3( Cell_4_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_6_io_out ),
       .io_nbrs_6( Cell_12_io_out ),
       .io_nbrs_7( Cell_13_io_out ),
       .io_nbrs_8( Cell_14_io_out ),
       .io_out( Cell_5_io_out )
  );
  Cell_1 Cell_6(.clk(clk),
       .io_in( T344 ),
       .io_in_val( T342 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( 1'h0 ),
       .io_nbrs_3( Cell_5_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_7_io_out ),
       .io_nbrs_6( Cell_13_io_out ),
       .io_nbrs_7( Cell_14_io_out ),
       .io_nbrs_8( Cell_15_io_out ),
       .io_out( Cell_6_io_out )
  );
  Cell_2 Cell_7(.clk(clk),
       .io_in( T338 ),
       .io_in_val( T336 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( 1'h0 ),
       .io_nbrs_2( Cell_0_io_out ),
       .io_nbrs_3( Cell_6_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_8_io_out ),
       .io_nbrs_6( Cell_14_io_out ),
       .io_nbrs_7( Cell_15_io_out ),
       .io_nbrs_8( Cell_16_io_out ),
       .io_out( Cell_7_io_out )
  );
  Cell_3 Cell_8(.clk(clk),
       .io_in( T332 ),
       .io_in_val( T330 ),
       .io_nbrs_0( 1'h0 ),
       .io_nbrs_1( Cell_0_io_out ),
       .io_nbrs_2( Cell_1_io_out ),
       .io_nbrs_3( Cell_7_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_9_io_out ),
       .io_nbrs_6( Cell_15_io_out ),
       .io_nbrs_7( Cell_16_io_out ),
       .io_nbrs_8( Cell_17_io_out ),
       .io_out( Cell_8_io_out )
  );
  Cell_4 Cell_9(.clk(clk),
       .io_in( T326 ),
       .io_in_val( T324 ),
       .io_nbrs_0( Cell_0_io_out ),
       .io_nbrs_1( Cell_1_io_out ),
       .io_nbrs_2( Cell_2_io_out ),
       .io_nbrs_3( Cell_8_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_10_io_out ),
       .io_nbrs_6( Cell_16_io_out ),
       .io_nbrs_7( Cell_17_io_out ),
       .io_nbrs_8( Cell_18_io_out ),
       .io_out( Cell_9_io_out )
  );
  Cell_4 Cell_10(.clk(clk),
       .io_in( T320 ),
       .io_in_val( T318 ),
       .io_nbrs_0( Cell_1_io_out ),
       .io_nbrs_1( Cell_2_io_out ),
       .io_nbrs_2( Cell_3_io_out ),
       .io_nbrs_3( Cell_9_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_11_io_out ),
       .io_nbrs_6( Cell_17_io_out ),
       .io_nbrs_7( Cell_18_io_out ),
       .io_nbrs_8( Cell_19_io_out ),
       .io_out( Cell_10_io_out )
  );
  Cell_4 Cell_11(.clk(clk),
       .io_in( T314 ),
       .io_in_val( T312 ),
       .io_nbrs_0( Cell_2_io_out ),
       .io_nbrs_1( Cell_3_io_out ),
       .io_nbrs_2( Cell_4_io_out ),
       .io_nbrs_3( Cell_10_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_12_io_out ),
       .io_nbrs_6( Cell_18_io_out ),
       .io_nbrs_7( Cell_19_io_out ),
       .io_nbrs_8( Cell_20_io_out ),
       .io_out( Cell_11_io_out )
  );
  Cell_4 Cell_12(.clk(clk),
       .io_in( T308 ),
       .io_in_val( T306 ),
       .io_nbrs_0( Cell_3_io_out ),
       .io_nbrs_1( Cell_4_io_out ),
       .io_nbrs_2( Cell_5_io_out ),
       .io_nbrs_3( Cell_11_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_13_io_out ),
       .io_nbrs_6( Cell_19_io_out ),
       .io_nbrs_7( Cell_20_io_out ),
       .io_nbrs_8( Cell_21_io_out ),
       .io_out( Cell_12_io_out )
  );
  Cell_4 Cell_13(.clk(clk),
       .io_in( T302 ),
       .io_in_val( T300 ),
       .io_nbrs_0( Cell_4_io_out ),
       .io_nbrs_1( Cell_5_io_out ),
       .io_nbrs_2( Cell_6_io_out ),
       .io_nbrs_3( Cell_12_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_14_io_out ),
       .io_nbrs_6( Cell_20_io_out ),
       .io_nbrs_7( Cell_21_io_out ),
       .io_nbrs_8( Cell_22_io_out ),
       .io_out( Cell_13_io_out )
  );
  Cell_4 Cell_14(.clk(clk),
       .io_in( T296 ),
       .io_in_val( T294 ),
       .io_nbrs_0( Cell_5_io_out ),
       .io_nbrs_1( Cell_6_io_out ),
       .io_nbrs_2( Cell_7_io_out ),
       .io_nbrs_3( Cell_13_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_15_io_out ),
       .io_nbrs_6( Cell_21_io_out ),
       .io_nbrs_7( Cell_22_io_out ),
       .io_nbrs_8( Cell_23_io_out ),
       .io_out( Cell_14_io_out )
  );
  Cell_4 Cell_15(.clk(clk),
       .io_in( T290 ),
       .io_in_val( T288 ),
       .io_nbrs_0( Cell_6_io_out ),
       .io_nbrs_1( Cell_7_io_out ),
       .io_nbrs_2( Cell_8_io_out ),
       .io_nbrs_3( Cell_14_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_16_io_out ),
       .io_nbrs_6( Cell_22_io_out ),
       .io_nbrs_7( Cell_23_io_out ),
       .io_nbrs_8( Cell_24_io_out ),
       .io_out( Cell_15_io_out )
  );
  Cell_4 Cell_16(.clk(clk),
       .io_in( T284 ),
       .io_in_val( T282 ),
       .io_nbrs_0( Cell_7_io_out ),
       .io_nbrs_1( Cell_8_io_out ),
       .io_nbrs_2( Cell_9_io_out ),
       .io_nbrs_3( Cell_15_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_17_io_out ),
       .io_nbrs_6( Cell_23_io_out ),
       .io_nbrs_7( Cell_24_io_out ),
       .io_nbrs_8( Cell_25_io_out ),
       .io_out( Cell_16_io_out )
  );
  Cell_4 Cell_17(.clk(clk),
       .io_in( T278 ),
       .io_in_val( T276 ),
       .io_nbrs_0( Cell_8_io_out ),
       .io_nbrs_1( Cell_9_io_out ),
       .io_nbrs_2( Cell_10_io_out ),
       .io_nbrs_3( Cell_16_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_18_io_out ),
       .io_nbrs_6( Cell_24_io_out ),
       .io_nbrs_7( Cell_25_io_out ),
       .io_nbrs_8( Cell_26_io_out ),
       .io_out( Cell_17_io_out )
  );
  Cell_4 Cell_18(.clk(clk),
       .io_in( T272 ),
       .io_in_val( T270 ),
       .io_nbrs_0( Cell_9_io_out ),
       .io_nbrs_1( Cell_10_io_out ),
       .io_nbrs_2( Cell_11_io_out ),
       .io_nbrs_3( Cell_17_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_19_io_out ),
       .io_nbrs_6( Cell_25_io_out ),
       .io_nbrs_7( Cell_26_io_out ),
       .io_nbrs_8( Cell_27_io_out ),
       .io_out( Cell_18_io_out )
  );
  Cell_4 Cell_19(.clk(clk),
       .io_in( T266 ),
       .io_in_val( T264 ),
       .io_nbrs_0( Cell_10_io_out ),
       .io_nbrs_1( Cell_11_io_out ),
       .io_nbrs_2( Cell_12_io_out ),
       .io_nbrs_3( Cell_18_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_20_io_out ),
       .io_nbrs_6( Cell_26_io_out ),
       .io_nbrs_7( Cell_27_io_out ),
       .io_nbrs_8( Cell_28_io_out ),
       .io_out( Cell_19_io_out )
  );
  Cell_4 Cell_20(.clk(clk),
       .io_in( T260 ),
       .io_in_val( T258 ),
       .io_nbrs_0( Cell_11_io_out ),
       .io_nbrs_1( Cell_12_io_out ),
       .io_nbrs_2( Cell_13_io_out ),
       .io_nbrs_3( Cell_19_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_21_io_out ),
       .io_nbrs_6( Cell_27_io_out ),
       .io_nbrs_7( Cell_28_io_out ),
       .io_nbrs_8( Cell_29_io_out ),
       .io_out( Cell_20_io_out )
  );
  Cell_4 Cell_21(.clk(clk),
       .io_in( T254 ),
       .io_in_val( T252 ),
       .io_nbrs_0( Cell_12_io_out ),
       .io_nbrs_1( Cell_13_io_out ),
       .io_nbrs_2( Cell_14_io_out ),
       .io_nbrs_3( Cell_20_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_22_io_out ),
       .io_nbrs_6( Cell_28_io_out ),
       .io_nbrs_7( Cell_29_io_out ),
       .io_nbrs_8( Cell_30_io_out ),
       .io_out( Cell_21_io_out )
  );
  Cell_4 Cell_22(.clk(clk),
       .io_in( T248 ),
       .io_in_val( T246 ),
       .io_nbrs_0( Cell_13_io_out ),
       .io_nbrs_1( Cell_14_io_out ),
       .io_nbrs_2( Cell_15_io_out ),
       .io_nbrs_3( Cell_21_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_23_io_out ),
       .io_nbrs_6( Cell_29_io_out ),
       .io_nbrs_7( Cell_30_io_out ),
       .io_nbrs_8( Cell_31_io_out ),
       .io_out( Cell_22_io_out )
  );
  Cell_4 Cell_23(.clk(clk),
       .io_in( T242 ),
       .io_in_val( T240 ),
       .io_nbrs_0( Cell_14_io_out ),
       .io_nbrs_1( Cell_15_io_out ),
       .io_nbrs_2( Cell_16_io_out ),
       .io_nbrs_3( Cell_22_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_24_io_out ),
       .io_nbrs_6( Cell_30_io_out ),
       .io_nbrs_7( Cell_31_io_out ),
       .io_nbrs_8( Cell_32_io_out ),
       .io_out( Cell_23_io_out )
  );
  Cell_4 Cell_24(.clk(clk),
       .io_in( T236 ),
       .io_in_val( T234 ),
       .io_nbrs_0( Cell_15_io_out ),
       .io_nbrs_1( Cell_16_io_out ),
       .io_nbrs_2( Cell_17_io_out ),
       .io_nbrs_3( Cell_23_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_25_io_out ),
       .io_nbrs_6( Cell_31_io_out ),
       .io_nbrs_7( Cell_32_io_out ),
       .io_nbrs_8( Cell_33_io_out ),
       .io_out( Cell_24_io_out )
  );
  Cell_4 Cell_25(.clk(clk),
       .io_in( T230 ),
       .io_in_val( T228 ),
       .io_nbrs_0( Cell_16_io_out ),
       .io_nbrs_1( Cell_17_io_out ),
       .io_nbrs_2( Cell_18_io_out ),
       .io_nbrs_3( Cell_24_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_26_io_out ),
       .io_nbrs_6( Cell_32_io_out ),
       .io_nbrs_7( Cell_33_io_out ),
       .io_nbrs_8( Cell_34_io_out ),
       .io_out( Cell_25_io_out )
  );
  Cell_4 Cell_26(.clk(clk),
       .io_in( T224 ),
       .io_in_val( T222 ),
       .io_nbrs_0( Cell_17_io_out ),
       .io_nbrs_1( Cell_18_io_out ),
       .io_nbrs_2( Cell_19_io_out ),
       .io_nbrs_3( Cell_25_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_27_io_out ),
       .io_nbrs_6( Cell_33_io_out ),
       .io_nbrs_7( Cell_34_io_out ),
       .io_nbrs_8( Cell_35_io_out ),
       .io_out( Cell_26_io_out )
  );
  Cell_4 Cell_27(.clk(clk),
       .io_in( T218 ),
       .io_in_val( T216 ),
       .io_nbrs_0( Cell_18_io_out ),
       .io_nbrs_1( Cell_19_io_out ),
       .io_nbrs_2( Cell_20_io_out ),
       .io_nbrs_3( Cell_26_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_28_io_out ),
       .io_nbrs_6( Cell_34_io_out ),
       .io_nbrs_7( Cell_35_io_out ),
       .io_nbrs_8( Cell_36_io_out ),
       .io_out( Cell_27_io_out )
  );
  Cell_4 Cell_28(.clk(clk),
       .io_in( T212 ),
       .io_in_val( T210 ),
       .io_nbrs_0( Cell_19_io_out ),
       .io_nbrs_1( Cell_20_io_out ),
       .io_nbrs_2( Cell_21_io_out ),
       .io_nbrs_3( Cell_27_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_29_io_out ),
       .io_nbrs_6( Cell_35_io_out ),
       .io_nbrs_7( Cell_36_io_out ),
       .io_nbrs_8( Cell_37_io_out ),
       .io_out( Cell_28_io_out )
  );
  Cell_4 Cell_29(.clk(clk),
       .io_in( T206 ),
       .io_in_val( T204 ),
       .io_nbrs_0( Cell_20_io_out ),
       .io_nbrs_1( Cell_21_io_out ),
       .io_nbrs_2( Cell_22_io_out ),
       .io_nbrs_3( Cell_28_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_30_io_out ),
       .io_nbrs_6( Cell_36_io_out ),
       .io_nbrs_7( Cell_37_io_out ),
       .io_nbrs_8( Cell_38_io_out ),
       .io_out( Cell_29_io_out )
  );
  Cell_4 Cell_30(.clk(clk),
       .io_in( T200 ),
       .io_in_val( T198 ),
       .io_nbrs_0( Cell_21_io_out ),
       .io_nbrs_1( Cell_22_io_out ),
       .io_nbrs_2( Cell_23_io_out ),
       .io_nbrs_3( Cell_29_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_31_io_out ),
       .io_nbrs_6( Cell_37_io_out ),
       .io_nbrs_7( Cell_38_io_out ),
       .io_nbrs_8( Cell_39_io_out ),
       .io_out( Cell_30_io_out )
  );
  Cell_4 Cell_31(.clk(clk),
       .io_in( T194 ),
       .io_in_val( T192 ),
       .io_nbrs_0( Cell_22_io_out ),
       .io_nbrs_1( Cell_23_io_out ),
       .io_nbrs_2( Cell_24_io_out ),
       .io_nbrs_3( Cell_30_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_32_io_out ),
       .io_nbrs_6( Cell_38_io_out ),
       .io_nbrs_7( Cell_39_io_out ),
       .io_nbrs_8( Cell_40_io_out ),
       .io_out( Cell_31_io_out )
  );
  Cell_4 Cell_32(.clk(clk),
       .io_in( T188 ),
       .io_in_val( T186 ),
       .io_nbrs_0( Cell_23_io_out ),
       .io_nbrs_1( Cell_24_io_out ),
       .io_nbrs_2( Cell_25_io_out ),
       .io_nbrs_3( Cell_31_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_33_io_out ),
       .io_nbrs_6( Cell_39_io_out ),
       .io_nbrs_7( Cell_40_io_out ),
       .io_nbrs_8( Cell_41_io_out ),
       .io_out( Cell_32_io_out )
  );
  Cell_4 Cell_33(.clk(clk),
       .io_in( T182 ),
       .io_in_val( T180 ),
       .io_nbrs_0( Cell_24_io_out ),
       .io_nbrs_1( Cell_25_io_out ),
       .io_nbrs_2( Cell_26_io_out ),
       .io_nbrs_3( Cell_32_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_34_io_out ),
       .io_nbrs_6( Cell_40_io_out ),
       .io_nbrs_7( Cell_41_io_out ),
       .io_nbrs_8( Cell_42_io_out ),
       .io_out( Cell_33_io_out )
  );
  Cell_4 Cell_34(.clk(clk),
       .io_in( T176 ),
       .io_in_val( T174 ),
       .io_nbrs_0( Cell_25_io_out ),
       .io_nbrs_1( Cell_26_io_out ),
       .io_nbrs_2( Cell_27_io_out ),
       .io_nbrs_3( Cell_33_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_35_io_out ),
       .io_nbrs_6( Cell_41_io_out ),
       .io_nbrs_7( Cell_42_io_out ),
       .io_nbrs_8( Cell_43_io_out ),
       .io_out( Cell_34_io_out )
  );
  Cell_4 Cell_35(.clk(clk),
       .io_in( T170 ),
       .io_in_val( T168 ),
       .io_nbrs_0( Cell_26_io_out ),
       .io_nbrs_1( Cell_27_io_out ),
       .io_nbrs_2( Cell_28_io_out ),
       .io_nbrs_3( Cell_34_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_36_io_out ),
       .io_nbrs_6( Cell_42_io_out ),
       .io_nbrs_7( Cell_43_io_out ),
       .io_nbrs_8( Cell_44_io_out ),
       .io_out( Cell_35_io_out )
  );
  Cell_4 Cell_36(.clk(clk),
       .io_in( T164 ),
       .io_in_val( T162 ),
       .io_nbrs_0( Cell_27_io_out ),
       .io_nbrs_1( Cell_28_io_out ),
       .io_nbrs_2( Cell_29_io_out ),
       .io_nbrs_3( Cell_35_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_37_io_out ),
       .io_nbrs_6( Cell_43_io_out ),
       .io_nbrs_7( Cell_44_io_out ),
       .io_nbrs_8( Cell_45_io_out ),
       .io_out( Cell_36_io_out )
  );
  Cell_4 Cell_37(.clk(clk),
       .io_in( T158 ),
       .io_in_val( T156 ),
       .io_nbrs_0( Cell_28_io_out ),
       .io_nbrs_1( Cell_29_io_out ),
       .io_nbrs_2( Cell_30_io_out ),
       .io_nbrs_3( Cell_36_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_38_io_out ),
       .io_nbrs_6( Cell_44_io_out ),
       .io_nbrs_7( Cell_45_io_out ),
       .io_nbrs_8( Cell_46_io_out ),
       .io_out( Cell_37_io_out )
  );
  Cell_4 Cell_38(.clk(clk),
       .io_in( T152 ),
       .io_in_val( T150 ),
       .io_nbrs_0( Cell_29_io_out ),
       .io_nbrs_1( Cell_30_io_out ),
       .io_nbrs_2( Cell_31_io_out ),
       .io_nbrs_3( Cell_37_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_39_io_out ),
       .io_nbrs_6( Cell_45_io_out ),
       .io_nbrs_7( Cell_46_io_out ),
       .io_nbrs_8( Cell_47_io_out ),
       .io_out( Cell_38_io_out )
  );
  Cell_4 Cell_39(.clk(clk),
       .io_in( T146 ),
       .io_in_val( T144 ),
       .io_nbrs_0( Cell_30_io_out ),
       .io_nbrs_1( Cell_31_io_out ),
       .io_nbrs_2( Cell_32_io_out ),
       .io_nbrs_3( Cell_38_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_40_io_out ),
       .io_nbrs_6( Cell_46_io_out ),
       .io_nbrs_7( Cell_47_io_out ),
       .io_nbrs_8( Cell_48_io_out ),
       .io_out( Cell_39_io_out )
  );
  Cell_4 Cell_40(.clk(clk),
       .io_in( T140 ),
       .io_in_val( T138 ),
       .io_nbrs_0( Cell_31_io_out ),
       .io_nbrs_1( Cell_32_io_out ),
       .io_nbrs_2( Cell_33_io_out ),
       .io_nbrs_3( Cell_39_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_41_io_out ),
       .io_nbrs_6( Cell_47_io_out ),
       .io_nbrs_7( Cell_48_io_out ),
       .io_nbrs_8( Cell_49_io_out ),
       .io_out( Cell_40_io_out )
  );
  Cell_4 Cell_41(.clk(clk),
       .io_in( T134 ),
       .io_in_val( T132 ),
       .io_nbrs_0( Cell_32_io_out ),
       .io_nbrs_1( Cell_33_io_out ),
       .io_nbrs_2( Cell_34_io_out ),
       .io_nbrs_3( Cell_40_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_42_io_out ),
       .io_nbrs_6( Cell_48_io_out ),
       .io_nbrs_7( Cell_49_io_out ),
       .io_nbrs_8( Cell_50_io_out ),
       .io_out( Cell_41_io_out )
  );
  Cell_4 Cell_42(.clk(clk),
       .io_in( T128 ),
       .io_in_val( T126 ),
       .io_nbrs_0( Cell_33_io_out ),
       .io_nbrs_1( Cell_34_io_out ),
       .io_nbrs_2( Cell_35_io_out ),
       .io_nbrs_3( Cell_41_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_43_io_out ),
       .io_nbrs_6( Cell_49_io_out ),
       .io_nbrs_7( Cell_50_io_out ),
       .io_nbrs_8( Cell_51_io_out ),
       .io_out( Cell_42_io_out )
  );
  Cell_4 Cell_43(.clk(clk),
       .io_in( T122 ),
       .io_in_val( T120 ),
       .io_nbrs_0( Cell_34_io_out ),
       .io_nbrs_1( Cell_35_io_out ),
       .io_nbrs_2( Cell_36_io_out ),
       .io_nbrs_3( Cell_42_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_44_io_out ),
       .io_nbrs_6( Cell_50_io_out ),
       .io_nbrs_7( Cell_51_io_out ),
       .io_nbrs_8( Cell_52_io_out ),
       .io_out( Cell_43_io_out )
  );
  Cell_4 Cell_44(.clk(clk),
       .io_in( T116 ),
       .io_in_val( T114 ),
       .io_nbrs_0( Cell_35_io_out ),
       .io_nbrs_1( Cell_36_io_out ),
       .io_nbrs_2( Cell_37_io_out ),
       .io_nbrs_3( Cell_43_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_45_io_out ),
       .io_nbrs_6( Cell_51_io_out ),
       .io_nbrs_7( Cell_52_io_out ),
       .io_nbrs_8( Cell_53_io_out ),
       .io_out( Cell_44_io_out )
  );
  Cell_4 Cell_45(.clk(clk),
       .io_in( T110 ),
       .io_in_val( T108 ),
       .io_nbrs_0( Cell_36_io_out ),
       .io_nbrs_1( Cell_37_io_out ),
       .io_nbrs_2( Cell_38_io_out ),
       .io_nbrs_3( Cell_44_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_46_io_out ),
       .io_nbrs_6( Cell_52_io_out ),
       .io_nbrs_7( Cell_53_io_out ),
       .io_nbrs_8( Cell_54_io_out ),
       .io_out( Cell_45_io_out )
  );
  Cell_4 Cell_46(.clk(clk),
       .io_in( T104 ),
       .io_in_val( T102 ),
       .io_nbrs_0( Cell_37_io_out ),
       .io_nbrs_1( Cell_38_io_out ),
       .io_nbrs_2( Cell_39_io_out ),
       .io_nbrs_3( Cell_45_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_47_io_out ),
       .io_nbrs_6( Cell_53_io_out ),
       .io_nbrs_7( Cell_54_io_out ),
       .io_nbrs_8( Cell_55_io_out ),
       .io_out( Cell_46_io_out )
  );
  Cell_4 Cell_47(.clk(clk),
       .io_in( T98 ),
       .io_in_val( T96 ),
       .io_nbrs_0( Cell_38_io_out ),
       .io_nbrs_1( Cell_39_io_out ),
       .io_nbrs_2( Cell_40_io_out ),
       .io_nbrs_3( Cell_46_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_48_io_out ),
       .io_nbrs_6( Cell_54_io_out ),
       .io_nbrs_7( Cell_55_io_out ),
       .io_nbrs_8( Cell_56_io_out ),
       .io_out( Cell_47_io_out )
  );
  Cell_4 Cell_48(.clk(clk),
       .io_in( T92 ),
       .io_in_val( T90 ),
       .io_nbrs_0( Cell_39_io_out ),
       .io_nbrs_1( Cell_40_io_out ),
       .io_nbrs_2( Cell_41_io_out ),
       .io_nbrs_3( Cell_47_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_49_io_out ),
       .io_nbrs_6( Cell_55_io_out ),
       .io_nbrs_7( Cell_56_io_out ),
       .io_nbrs_8( Cell_57_io_out ),
       .io_out( Cell_48_io_out )
  );
  Cell_4 Cell_49(.clk(clk),
       .io_in( T86 ),
       .io_in_val( T84 ),
       .io_nbrs_0( Cell_40_io_out ),
       .io_nbrs_1( Cell_41_io_out ),
       .io_nbrs_2( Cell_42_io_out ),
       .io_nbrs_3( Cell_48_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_50_io_out ),
       .io_nbrs_6( Cell_56_io_out ),
       .io_nbrs_7( Cell_57_io_out ),
       .io_nbrs_8( Cell_58_io_out ),
       .io_out( Cell_49_io_out )
  );
  Cell_4 Cell_50(.clk(clk),
       .io_in( T80 ),
       .io_in_val( T78 ),
       .io_nbrs_0( Cell_41_io_out ),
       .io_nbrs_1( Cell_42_io_out ),
       .io_nbrs_2( Cell_43_io_out ),
       .io_nbrs_3( Cell_49_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_51_io_out ),
       .io_nbrs_6( Cell_57_io_out ),
       .io_nbrs_7( Cell_58_io_out ),
       .io_nbrs_8( Cell_59_io_out ),
       .io_out( Cell_50_io_out )
  );
  Cell_4 Cell_51(.clk(clk),
       .io_in( T74 ),
       .io_in_val( T72 ),
       .io_nbrs_0( Cell_42_io_out ),
       .io_nbrs_1( Cell_43_io_out ),
       .io_nbrs_2( Cell_44_io_out ),
       .io_nbrs_3( Cell_50_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_52_io_out ),
       .io_nbrs_6( Cell_58_io_out ),
       .io_nbrs_7( Cell_59_io_out ),
       .io_nbrs_8( Cell_60_io_out ),
       .io_out( Cell_51_io_out )
  );
  Cell_4 Cell_52(.clk(clk),
       .io_in( T68 ),
       .io_in_val( T66 ),
       .io_nbrs_0( Cell_43_io_out ),
       .io_nbrs_1( Cell_44_io_out ),
       .io_nbrs_2( Cell_45_io_out ),
       .io_nbrs_3( Cell_51_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_53_io_out ),
       .io_nbrs_6( Cell_59_io_out ),
       .io_nbrs_7( Cell_60_io_out ),
       .io_nbrs_8( Cell_61_io_out ),
       .io_out( Cell_52_io_out )
  );
  Cell_4 Cell_53(.clk(clk),
       .io_in( T62 ),
       .io_in_val( T60 ),
       .io_nbrs_0( Cell_44_io_out ),
       .io_nbrs_1( Cell_45_io_out ),
       .io_nbrs_2( Cell_46_io_out ),
       .io_nbrs_3( Cell_52_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_54_io_out ),
       .io_nbrs_6( Cell_60_io_out ),
       .io_nbrs_7( Cell_61_io_out ),
       .io_nbrs_8( Cell_62_io_out ),
       .io_out( Cell_53_io_out )
  );
  Cell_4 Cell_54(.clk(clk),
       .io_in( T56 ),
       .io_in_val( T54 ),
       .io_nbrs_0( Cell_45_io_out ),
       .io_nbrs_1( Cell_46_io_out ),
       .io_nbrs_2( Cell_47_io_out ),
       .io_nbrs_3( Cell_53_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_55_io_out ),
       .io_nbrs_6( Cell_61_io_out ),
       .io_nbrs_7( Cell_62_io_out ),
       .io_nbrs_8( Cell_63_io_out ),
       .io_out( Cell_54_io_out )
  );
  Cell_5 Cell_55(.clk(clk),
       .io_in( T50 ),
       .io_in_val( T48 ),
       .io_nbrs_0( Cell_46_io_out ),
       .io_nbrs_1( Cell_47_io_out ),
       .io_nbrs_2( Cell_48_io_out ),
       .io_nbrs_3( Cell_54_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_56_io_out ),
       .io_nbrs_6( Cell_62_io_out ),
       .io_nbrs_7( Cell_63_io_out ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_55_io_out )
  );
  Cell_6 Cell_56(.clk(clk),
       .io_in( T44 ),
       .io_in_val( T42 ),
       .io_nbrs_0( Cell_47_io_out ),
       .io_nbrs_1( Cell_48_io_out ),
       .io_nbrs_2( Cell_49_io_out ),
       .io_nbrs_3( Cell_55_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_57_io_out ),
       .io_nbrs_6( Cell_63_io_out ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_56_io_out )
  );
  Cell_7 Cell_57(.clk(clk),
       .io_in( T38 ),
       .io_in_val( T36 ),
       .io_nbrs_0( Cell_48_io_out ),
       .io_nbrs_1( Cell_49_io_out ),
       .io_nbrs_2( Cell_50_io_out ),
       .io_nbrs_3( Cell_56_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_58_io_out ),
       .io_nbrs_6( 1'h0 ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_57_io_out )
  );
  Cell_7 Cell_58(.clk(clk),
       .io_in( T32 ),
       .io_in_val( T30 ),
       .io_nbrs_0( Cell_49_io_out ),
       .io_nbrs_1( Cell_50_io_out ),
       .io_nbrs_2( Cell_51_io_out ),
       .io_nbrs_3( Cell_57_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_59_io_out ),
       .io_nbrs_6( 1'h0 ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_58_io_out )
  );
  Cell_7 Cell_59(.clk(clk),
       .io_in( T26 ),
       .io_in_val( T24 ),
       .io_nbrs_0( Cell_50_io_out ),
       .io_nbrs_1( Cell_51_io_out ),
       .io_nbrs_2( Cell_52_io_out ),
       .io_nbrs_3( Cell_58_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_60_io_out ),
       .io_nbrs_6( 1'h0 ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_59_io_out )
  );
  Cell_7 Cell_60(.clk(clk),
       .io_in( T20 ),
       .io_in_val( T18 ),
       .io_nbrs_0( Cell_51_io_out ),
       .io_nbrs_1( Cell_52_io_out ),
       .io_nbrs_2( Cell_53_io_out ),
       .io_nbrs_3( Cell_59_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_61_io_out ),
       .io_nbrs_6( 1'h0 ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_60_io_out )
  );
  Cell_7 Cell_61(.clk(clk),
       .io_in( T14 ),
       .io_in_val( T12 ),
       .io_nbrs_0( Cell_52_io_out ),
       .io_nbrs_1( Cell_53_io_out ),
       .io_nbrs_2( Cell_54_io_out ),
       .io_nbrs_3( Cell_60_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_62_io_out ),
       .io_nbrs_6( 1'h0 ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_61_io_out )
  );
  Cell_7 Cell_62(.clk(clk),
       .io_in( T8 ),
       .io_in_val( T6 ),
       .io_nbrs_0( Cell_53_io_out ),
       .io_nbrs_1( Cell_54_io_out ),
       .io_nbrs_2( Cell_55_io_out ),
       .io_nbrs_3( Cell_61_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( Cell_63_io_out ),
       .io_nbrs_6( 1'h0 ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_62_io_out )
  );
  Cell_8 Cell_63(.clk(clk),
       .io_in( T2 ),
       .io_in_val( T0 ),
       .io_nbrs_0( Cell_54_io_out ),
       .io_nbrs_1( Cell_55_io_out ),
       .io_nbrs_2( Cell_56_io_out ),
       .io_nbrs_3( Cell_62_io_out ),
       .io_nbrs_4( 1'h0 ),
       .io_nbrs_5( 1'h0 ),
       .io_nbrs_6( 1'h0 ),
       .io_nbrs_7( 1'h0 ),
       .io_nbrs_8( 1'h0 ),
       .io_out( Cell_63_io_out )
  );

  always @(posedge clk) begin
    R387 <= reset ? 5'h0 : T388;
    if(reset) begin
      check_out <= 64'h1;
    end else if(T392) begin
      check_out <= T394;
    end
    if(reset) begin
      is_full <= 1'h0;
    end else if(T465) begin
      is_full <= T529;
    end
  end
endmodule

module Controller(input clk, input reset,
    input [63:0] io_rx_dat_int,
    input  io_rx_val,
    output[63:0] io_tx_dat_int,
    output io_tx_val
);

  wire T0;
  wire T1;
  wire Fifo_19_io_deq_val;
  wire Mapper_19_io_rx_rdy;
  wire T2;
  wire[63:0] Fifo_19_io_deq_dat_int;
  wire T3;
  wire T4;
  wire Fifo_18_io_deq_val;
  wire Mapper_18_io_rx_rdy;
  wire T5;
  wire[63:0] Fifo_18_io_deq_dat_int;
  wire T6;
  wire T7;
  wire Fifo_17_io_deq_val;
  wire Mapper_17_io_rx_rdy;
  wire T8;
  wire[63:0] Fifo_17_io_deq_dat_int;
  wire T9;
  wire T10;
  wire Fifo_16_io_deq_val;
  wire Mapper_16_io_rx_rdy;
  wire T11;
  wire[63:0] Fifo_16_io_deq_dat_int;
  wire T12;
  wire T13;
  wire Fifo_15_io_deq_val;
  wire Mapper_15_io_rx_rdy;
  wire T14;
  wire[63:0] Fifo_15_io_deq_dat_int;
  wire T15;
  wire T16;
  wire Fifo_14_io_deq_val;
  wire Mapper_14_io_rx_rdy;
  wire T17;
  wire[63:0] Fifo_14_io_deq_dat_int;
  wire T18;
  wire T19;
  wire Fifo_13_io_deq_val;
  wire Mapper_13_io_rx_rdy;
  wire T20;
  wire[63:0] Fifo_13_io_deq_dat_int;
  wire T21;
  wire T22;
  wire Fifo_12_io_deq_val;
  wire Mapper_12_io_rx_rdy;
  wire T23;
  wire[63:0] Fifo_12_io_deq_dat_int;
  wire T24;
  wire T25;
  wire Fifo_11_io_deq_val;
  wire Mapper_11_io_rx_rdy;
  wire T26;
  wire[63:0] Fifo_11_io_deq_dat_int;
  wire T27;
  wire T28;
  wire Fifo_10_io_deq_val;
  wire Mapper_10_io_rx_rdy;
  wire T29;
  wire[63:0] Fifo_10_io_deq_dat_int;
  wire T30;
  wire T31;
  wire Fifo_9_io_deq_val;
  wire Mapper_9_io_rx_rdy;
  wire T32;
  wire[63:0] Fifo_9_io_deq_dat_int;
  wire T33;
  wire T34;
  wire Fifo_8_io_deq_val;
  wire Mapper_8_io_rx_rdy;
  wire T35;
  wire[63:0] Fifo_8_io_deq_dat_int;
  wire T36;
  wire T37;
  wire Fifo_7_io_deq_val;
  wire Mapper_7_io_rx_rdy;
  wire T38;
  wire[63:0] Fifo_7_io_deq_dat_int;
  wire T39;
  wire T40;
  wire Fifo_6_io_deq_val;
  wire Mapper_6_io_rx_rdy;
  wire T41;
  wire[63:0] Fifo_6_io_deq_dat_int;
  wire T42;
  wire T43;
  wire Fifo_5_io_deq_val;
  wire Mapper_5_io_rx_rdy;
  wire T44;
  wire[63:0] Fifo_5_io_deq_dat_int;
  wire T45;
  wire T46;
  wire Fifo_4_io_deq_val;
  wire Mapper_4_io_rx_rdy;
  wire T47;
  wire[63:0] Fifo_4_io_deq_dat_int;
  wire T48;
  wire T49;
  wire Fifo_3_io_deq_val;
  wire Mapper_3_io_rx_rdy;
  wire T50;
  wire[63:0] Fifo_3_io_deq_dat_int;
  wire T51;
  wire T52;
  wire Fifo_2_io_deq_val;
  wire Mapper_2_io_rx_rdy;
  wire T53;
  wire[63:0] Fifo_2_io_deq_dat_int;
  wire T54;
  wire T55;
  wire Fifo_1_io_deq_val;
  wire Mapper_1_io_rx_rdy;
  wire T56;
  wire[63:0] Fifo_1_io_deq_dat_int;
  wire T57;
  wire T58;
  wire Fifo_0_io_deq_val;
  wire Mapper_0_io_rx_rdy;
  wire T59;
  wire[63:0] Fifo_0_io_deq_dat_int;
  wire[63:0] Mapper_19_io_tx_dat_int;
  wire T60;
  wire T61;
  wire Fifo_39_io_deq_val;
  wire T62;
  wire[4:0] index;
  wire[4:0] T63;
  wire[4:0] T64;
  wire[4:0] T65;
  wire[4:0] T66;
  wire[3:0] T67;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire[3:0] T74;
  wire[3:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire[1:0] T83;
  wire T84;
  wire f_out_deq_rdy_1;
  wire T85;
  wire Fifo_21_io_deq_val;
  wire T86;
  wire f_out_deq_rdy_2;
  wire T87;
  wire Fifo_22_io_deq_val;
  wire T88;
  wire f_out_deq_rdy_3;
  wire T89;
  wire Fifo_23_io_deq_val;
  wire T90;
  wire f_out_deq_rdy_4;
  wire T91;
  wire Fifo_24_io_deq_val;
  wire T92;
  wire f_out_deq_rdy_5;
  wire T93;
  wire Fifo_25_io_deq_val;
  wire T94;
  wire f_out_deq_rdy_6;
  wire T95;
  wire Fifo_26_io_deq_val;
  wire T96;
  wire f_out_deq_rdy_7;
  wire T97;
  wire Fifo_27_io_deq_val;
  wire T98;
  wire f_out_deq_rdy_8;
  wire T99;
  wire Fifo_28_io_deq_val;
  wire T100;
  wire f_out_deq_rdy_9;
  wire T101;
  wire Fifo_29_io_deq_val;
  wire T102;
  wire f_out_deq_rdy_10;
  wire T103;
  wire Fifo_30_io_deq_val;
  wire T104;
  wire f_out_deq_rdy_11;
  wire T105;
  wire Fifo_31_io_deq_val;
  wire T106;
  wire f_out_deq_rdy_12;
  wire T107;
  wire Fifo_32_io_deq_val;
  wire T108;
  wire f_out_deq_rdy_13;
  wire T109;
  wire Fifo_33_io_deq_val;
  wire T110;
  wire f_out_deq_rdy_14;
  wire T111;
  wire Fifo_34_io_deq_val;
  wire T112;
  wire f_out_deq_rdy_15;
  wire T113;
  wire Fifo_35_io_deq_val;
  wire T114;
  wire f_out_deq_rdy_16;
  wire T115;
  wire Fifo_36_io_deq_val;
  wire T116;
  wire f_out_deq_rdy_17;
  wire T117;
  wire Fifo_37_io_deq_val;
  wire T118;
  wire f_out_deq_rdy_18;
  wire T119;
  wire Fifo_38_io_deq_val;
  wire T120;
  wire f_out_deq_rdy_19;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire Fifo_39_io_enq_rdy;
  wire Mapper_19_io_tx_val;
  wire T125;
  wire[63:0] Mapper_18_io_tx_dat_int;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire Fifo_38_io_enq_rdy;
  wire Mapper_18_io_tx_val;
  wire T132;
  wire[63:0] Mapper_17_io_tx_dat_int;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire Fifo_37_io_enq_rdy;
  wire Mapper_17_io_tx_val;
  wire T139;
  wire[63:0] Mapper_16_io_tx_dat_int;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire Fifo_36_io_enq_rdy;
  wire Mapper_16_io_tx_val;
  wire T146;
  wire[63:0] Mapper_15_io_tx_dat_int;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire Fifo_35_io_enq_rdy;
  wire Mapper_15_io_tx_val;
  wire T153;
  wire[63:0] Mapper_14_io_tx_dat_int;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire Fifo_34_io_enq_rdy;
  wire Mapper_14_io_tx_val;
  wire T160;
  wire[63:0] Mapper_13_io_tx_dat_int;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire Fifo_33_io_enq_rdy;
  wire Mapper_13_io_tx_val;
  wire T167;
  wire[63:0] Mapper_12_io_tx_dat_int;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire Fifo_32_io_enq_rdy;
  wire Mapper_12_io_tx_val;
  wire T174;
  wire[63:0] Mapper_11_io_tx_dat_int;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire Fifo_31_io_enq_rdy;
  wire Mapper_11_io_tx_val;
  wire T181;
  wire[63:0] Mapper_10_io_tx_dat_int;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire Fifo_30_io_enq_rdy;
  wire Mapper_10_io_tx_val;
  wire T188;
  wire[63:0] Mapper_9_io_tx_dat_int;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire Fifo_29_io_enq_rdy;
  wire Mapper_9_io_tx_val;
  wire T195;
  wire[63:0] Mapper_8_io_tx_dat_int;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire Fifo_28_io_enq_rdy;
  wire Mapper_8_io_tx_val;
  wire T202;
  wire[63:0] Mapper_7_io_tx_dat_int;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire Fifo_27_io_enq_rdy;
  wire Mapper_7_io_tx_val;
  wire T209;
  wire[63:0] Mapper_6_io_tx_dat_int;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire Fifo_26_io_enq_rdy;
  wire Mapper_6_io_tx_val;
  wire T216;
  wire[63:0] Mapper_5_io_tx_dat_int;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire Fifo_25_io_enq_rdy;
  wire Mapper_5_io_tx_val;
  wire T223;
  wire[63:0] Mapper_4_io_tx_dat_int;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire Fifo_24_io_enq_rdy;
  wire Mapper_4_io_tx_val;
  wire T230;
  wire[63:0] Mapper_3_io_tx_dat_int;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire Fifo_23_io_enq_rdy;
  wire Mapper_3_io_tx_val;
  wire T237;
  wire[63:0] Mapper_2_io_tx_dat_int;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire Fifo_22_io_enq_rdy;
  wire Mapper_2_io_tx_val;
  wire T244;
  wire[63:0] Mapper_1_io_tx_dat_int;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire Fifo_21_io_enq_rdy;
  wire Mapper_1_io_tx_val;
  wire T251;
  wire[63:0] Mapper_0_io_tx_dat_int;
  wire T252;
  wire T253;
  wire Fifo_20_io_deq_val;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire Fifo_20_io_enq_rdy;
  wire Mapper_0_io_tx_val;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire Fifo_19_io_enq_rdy;
  wire T262;
  wire T263;
  reg[4:0] inCounter;
  wire T264;
  wire T265;
  wire T266;
  wire Fifo_18_io_enq_rdy;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire Fifo_17_io_enq_rdy;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire Fifo_16_io_enq_rdy;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire Fifo_15_io_enq_rdy;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire Fifo_14_io_enq_rdy;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire Fifo_13_io_enq_rdy;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire Fifo_12_io_enq_rdy;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire Fifo_11_io_enq_rdy;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire Fifo_10_io_enq_rdy;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire Fifo_9_io_enq_rdy;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire Fifo_8_io_enq_rdy;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire Fifo_7_io_enq_rdy;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire Fifo_6_io_enq_rdy;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire Fifo_5_io_enq_rdy;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire Fifo_4_io_enq_rdy;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire Fifo_3_io_enq_rdy;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire Fifo_2_io_enq_rdy;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire Fifo_1_io_enq_rdy;
  wire T335;
  wire T336;
  wire T337;
  wire Fifo_0_io_enq_rdy;
  wire T338;
  wire T339;
  wire[4:0] T340;
  wire[4:0] T341;
  wire[4:0] T342;
  wire[4:0] T343;
  wire[4:0] T344;
  wire[4:0] T345;
  wire[4:0] T346;
  wire[4:0] T347;
  wire[4:0] T348;
  wire[4:0] T349;
  wire[4:0] T350;
  wire[4:0] T351;
  wire[4:0] T352;
  wire[4:0] T353;
  wire[4:0] T354;
  wire[4:0] T355;
  wire[4:0] T356;
  wire[4:0] T357;
  wire[4:0] T358;
  wire[4:0] T359;
  wire[4:0] T360;
  wire T361;
  wire[4:0] T362;
  wire[4:0] T363;
  wire T364;
  wire[4:0] T365;
  wire[4:0] T366;
  wire T367;
  wire[4:0] T368;
  wire[4:0] T369;
  wire T370;
  wire[4:0] T371;
  wire[4:0] T372;
  wire T373;
  wire[4:0] T374;
  wire[4:0] T375;
  wire T376;
  wire[4:0] T377;
  wire[4:0] T378;
  wire T379;
  wire[4:0] T380;
  wire[4:0] T381;
  wire T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire T385;
  wire[4:0] T386;
  wire[4:0] T387;
  wire T388;
  wire[4:0] T389;
  wire[4:0] T390;
  wire T391;
  wire[4:0] T392;
  wire[4:0] T393;
  wire T394;
  wire[4:0] T395;
  wire[4:0] T396;
  wire T397;
  wire[4:0] T398;
  wire[4:0] T399;
  wire T400;
  wire[4:0] T401;
  wire[4:0] T402;
  wire T403;
  wire[4:0] T404;
  wire[4:0] T405;
  wire T406;
  wire[4:0] T407;
  wire[4:0] T408;
  wire T409;
  wire[4:0] T410;
  wire[4:0] T411;
  wire T412;
  wire[4:0] T413;
  wire[4:0] T414;
  wire T415;
  wire[4:0] T416;
  wire[4:0] T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire[63:0] T496;
  wire[63:0] T497;
  wire[63:0] T498;
  wire[63:0] T499;
  wire[63:0] T500;
  wire[63:0] T501;
  wire[63:0] T502;
  wire[63:0] T503;
  wire[63:0] T504;
  wire[63:0] T505;
  wire[63:0] T506;
  wire[63:0] T507;
  wire[63:0] T508;
  wire[63:0] T509;
  wire[63:0] T510;
  wire[63:0] T511;
  wire[63:0] T512;
  wire[63:0] T513;
  wire[63:0] T514;
  wire[63:0] T515;
  wire[63:0] Fifo_20_io_deq_dat_int;
  wire[63:0] Fifo_21_io_deq_dat_int;
  wire[63:0] Fifo_22_io_deq_dat_int;
  wire[63:0] Fifo_23_io_deq_dat_int;
  wire[63:0] Fifo_24_io_deq_dat_int;
  wire[63:0] Fifo_25_io_deq_dat_int;
  wire[63:0] Fifo_26_io_deq_dat_int;
  wire[63:0] Fifo_27_io_deq_dat_int;
  wire[63:0] Fifo_28_io_deq_dat_int;
  wire[63:0] Fifo_29_io_deq_dat_int;
  wire[63:0] Fifo_30_io_deq_dat_int;
  wire[63:0] Fifo_31_io_deq_dat_int;
  wire[63:0] Fifo_32_io_deq_dat_int;
  wire[63:0] Fifo_33_io_deq_dat_int;
  wire[63:0] Fifo_34_io_deq_dat_int;
  wire[63:0] Fifo_35_io_deq_dat_int;
  wire[63:0] Fifo_36_io_deq_dat_int;
  wire[63:0] Fifo_37_io_deq_dat_int;
  wire[63:0] Fifo_38_io_deq_dat_int;
  wire[63:0] Fifo_39_io_deq_dat_int;

  assign T0 = T2 ? 1'h0 : T1;
  assign T1 = Mapper_19_io_rx_rdy && Fifo_19_io_deq_val;
  assign T2 = ! T1;
  assign T3 = T5 ? 1'h0 : T4;
  assign T4 = Mapper_18_io_rx_rdy && Fifo_18_io_deq_val;
  assign T5 = ! T4;
  assign T6 = T8 ? 1'h0 : T7;
  assign T7 = Mapper_17_io_rx_rdy && Fifo_17_io_deq_val;
  assign T8 = ! T7;
  assign T9 = T11 ? 1'h0 : T10;
  assign T10 = Mapper_16_io_rx_rdy && Fifo_16_io_deq_val;
  assign T11 = ! T10;
  assign T12 = T14 ? 1'h0 : T13;
  assign T13 = Mapper_15_io_rx_rdy && Fifo_15_io_deq_val;
  assign T14 = ! T13;
  assign T15 = T17 ? 1'h0 : T16;
  assign T16 = Mapper_14_io_rx_rdy && Fifo_14_io_deq_val;
  assign T17 = ! T16;
  assign T18 = T20 ? 1'h0 : T19;
  assign T19 = Mapper_13_io_rx_rdy && Fifo_13_io_deq_val;
  assign T20 = ! T19;
  assign T21 = T23 ? 1'h0 : T22;
  assign T22 = Mapper_12_io_rx_rdy && Fifo_12_io_deq_val;
  assign T23 = ! T22;
  assign T24 = T26 ? 1'h0 : T25;
  assign T25 = Mapper_11_io_rx_rdy && Fifo_11_io_deq_val;
  assign T26 = ! T25;
  assign T27 = T29 ? 1'h0 : T28;
  assign T28 = Mapper_10_io_rx_rdy && Fifo_10_io_deq_val;
  assign T29 = ! T28;
  assign T30 = T32 ? 1'h0 : T31;
  assign T31 = Mapper_9_io_rx_rdy && Fifo_9_io_deq_val;
  assign T32 = ! T31;
  assign T33 = T35 ? 1'h0 : T34;
  assign T34 = Mapper_8_io_rx_rdy && Fifo_8_io_deq_val;
  assign T35 = ! T34;
  assign T36 = T38 ? 1'h0 : T37;
  assign T37 = Mapper_7_io_rx_rdy && Fifo_7_io_deq_val;
  assign T38 = ! T37;
  assign T39 = T41 ? 1'h0 : T40;
  assign T40 = Mapper_6_io_rx_rdy && Fifo_6_io_deq_val;
  assign T41 = ! T40;
  assign T42 = T44 ? 1'h0 : T43;
  assign T43 = Mapper_5_io_rx_rdy && Fifo_5_io_deq_val;
  assign T44 = ! T43;
  assign T45 = T47 ? 1'h0 : T46;
  assign T46 = Mapper_4_io_rx_rdy && Fifo_4_io_deq_val;
  assign T47 = ! T46;
  assign T48 = T50 ? 1'h0 : T49;
  assign T49 = Mapper_3_io_rx_rdy && Fifo_3_io_deq_val;
  assign T50 = ! T49;
  assign T51 = T53 ? 1'h0 : T52;
  assign T52 = Mapper_2_io_rx_rdy && Fifo_2_io_deq_val;
  assign T53 = ! T52;
  assign T54 = T56 ? 1'h0 : T55;
  assign T55 = Mapper_1_io_rx_rdy && Fifo_1_io_deq_val;
  assign T56 = ! T55;
  assign T57 = T59 ? 1'h0 : T58;
  assign T58 = Mapper_0_io_rx_rdy && Fifo_0_io_deq_val;
  assign T59 = ! T58;
  assign T60 = T122 ? 1'h0 : T61;
  assign T61 = T62 && Fifo_39_io_deq_val;
  assign T62 = 5'h13 == index;
  assign index = T120 ? 5'h13 : T63;
  assign T63 = T118 ? 5'h12 : T64;
  assign T64 = T116 ? 5'h11 : T65;
  assign T65 = T114 ? 5'h10 : T66;
  assign T66 = {1'h0, T67};
  assign T67 = T112 ? 4'hf : T68;
  assign T68 = T110 ? 4'he : T69;
  assign T69 = T108 ? 4'hd : T70;
  assign T70 = T106 ? 4'hc : T71;
  assign T71 = T104 ? 4'hb : T72;
  assign T72 = T102 ? 4'ha : T73;
  assign T73 = T100 ? 4'h9 : T74;
  assign T74 = T98 ? 4'h8 : T75;
  assign T75 = {1'h0, T76};
  assign T76 = T96 ? 3'h7 : T77;
  assign T77 = T94 ? 3'h6 : T78;
  assign T78 = T92 ? 3'h5 : T79;
  assign T79 = T90 ? 3'h4 : T80;
  assign T80 = {1'h0, T81};
  assign T81 = T88 ? 2'h3 : T82;
  assign T82 = T86 ? 2'h2 : T83;
  assign T83 = {1'h0, T84};
  assign T84 = f_out_deq_rdy_1 == 1'h1;
  assign f_out_deq_rdy_1 = T85;
  assign T85 = Fifo_21_io_deq_val;
  assign T86 = f_out_deq_rdy_2 == 1'h1;
  assign f_out_deq_rdy_2 = T87;
  assign T87 = Fifo_22_io_deq_val;
  assign T88 = f_out_deq_rdy_3 == 1'h1;
  assign f_out_deq_rdy_3 = T89;
  assign T89 = Fifo_23_io_deq_val;
  assign T90 = f_out_deq_rdy_4 == 1'h1;
  assign f_out_deq_rdy_4 = T91;
  assign T91 = Fifo_24_io_deq_val;
  assign T92 = f_out_deq_rdy_5 == 1'h1;
  assign f_out_deq_rdy_5 = T93;
  assign T93 = Fifo_25_io_deq_val;
  assign T94 = f_out_deq_rdy_6 == 1'h1;
  assign f_out_deq_rdy_6 = T95;
  assign T95 = Fifo_26_io_deq_val;
  assign T96 = f_out_deq_rdy_7 == 1'h1;
  assign f_out_deq_rdy_7 = T97;
  assign T97 = Fifo_27_io_deq_val;
  assign T98 = f_out_deq_rdy_8 == 1'h1;
  assign f_out_deq_rdy_8 = T99;
  assign T99 = Fifo_28_io_deq_val;
  assign T100 = f_out_deq_rdy_9 == 1'h1;
  assign f_out_deq_rdy_9 = T101;
  assign T101 = Fifo_29_io_deq_val;
  assign T102 = f_out_deq_rdy_10 == 1'h1;
  assign f_out_deq_rdy_10 = T103;
  assign T103 = Fifo_30_io_deq_val;
  assign T104 = f_out_deq_rdy_11 == 1'h1;
  assign f_out_deq_rdy_11 = T105;
  assign T105 = Fifo_31_io_deq_val;
  assign T106 = f_out_deq_rdy_12 == 1'h1;
  assign f_out_deq_rdy_12 = T107;
  assign T107 = Fifo_32_io_deq_val;
  assign T108 = f_out_deq_rdy_13 == 1'h1;
  assign f_out_deq_rdy_13 = T109;
  assign T109 = Fifo_33_io_deq_val;
  assign T110 = f_out_deq_rdy_14 == 1'h1;
  assign f_out_deq_rdy_14 = T111;
  assign T111 = Fifo_34_io_deq_val;
  assign T112 = f_out_deq_rdy_15 == 1'h1;
  assign f_out_deq_rdy_15 = T113;
  assign T113 = Fifo_35_io_deq_val;
  assign T114 = f_out_deq_rdy_16 == 1'h1;
  assign f_out_deq_rdy_16 = T115;
  assign T115 = Fifo_36_io_deq_val;
  assign T116 = f_out_deq_rdy_17 == 1'h1;
  assign f_out_deq_rdy_17 = T117;
  assign T117 = Fifo_37_io_deq_val;
  assign T118 = f_out_deq_rdy_18 == 1'h1;
  assign f_out_deq_rdy_18 = T119;
  assign T119 = Fifo_38_io_deq_val;
  assign T120 = f_out_deq_rdy_19 == 1'h1;
  assign f_out_deq_rdy_19 = T121;
  assign T121 = Fifo_39_io_deq_val;
  assign T122 = ! T61;
  assign T123 = T125 ? 1'h0 : T124;
  assign T124 = Mapper_19_io_tx_val && Fifo_39_io_enq_rdy;
  assign T125 = ! T124;
  assign T126 = T129 ? 1'h0 : T127;
  assign T127 = T128 && Fifo_38_io_deq_val;
  assign T128 = 5'h12 == index;
  assign T129 = ! T127;
  assign T130 = T132 ? 1'h0 : T131;
  assign T131 = Mapper_18_io_tx_val && Fifo_38_io_enq_rdy;
  assign T132 = ! T131;
  assign T133 = T136 ? 1'h0 : T134;
  assign T134 = T135 && Fifo_37_io_deq_val;
  assign T135 = 5'h11 == index;
  assign T136 = ! T134;
  assign T137 = T139 ? 1'h0 : T138;
  assign T138 = Mapper_17_io_tx_val && Fifo_37_io_enq_rdy;
  assign T139 = ! T138;
  assign T140 = T143 ? 1'h0 : T141;
  assign T141 = T142 && Fifo_36_io_deq_val;
  assign T142 = 5'h10 == index;
  assign T143 = ! T141;
  assign T144 = T146 ? 1'h0 : T145;
  assign T145 = Mapper_16_io_tx_val && Fifo_36_io_enq_rdy;
  assign T146 = ! T145;
  assign T147 = T150 ? 1'h0 : T148;
  assign T148 = T149 && Fifo_35_io_deq_val;
  assign T149 = 5'hf == index;
  assign T150 = ! T148;
  assign T151 = T153 ? 1'h0 : T152;
  assign T152 = Mapper_15_io_tx_val && Fifo_35_io_enq_rdy;
  assign T153 = ! T152;
  assign T154 = T157 ? 1'h0 : T155;
  assign T155 = T156 && Fifo_34_io_deq_val;
  assign T156 = 5'he == index;
  assign T157 = ! T155;
  assign T158 = T160 ? 1'h0 : T159;
  assign T159 = Mapper_14_io_tx_val && Fifo_34_io_enq_rdy;
  assign T160 = ! T159;
  assign T161 = T164 ? 1'h0 : T162;
  assign T162 = T163 && Fifo_33_io_deq_val;
  assign T163 = 5'hd == index;
  assign T164 = ! T162;
  assign T165 = T167 ? 1'h0 : T166;
  assign T166 = Mapper_13_io_tx_val && Fifo_33_io_enq_rdy;
  assign T167 = ! T166;
  assign T168 = T171 ? 1'h0 : T169;
  assign T169 = T170 && Fifo_32_io_deq_val;
  assign T170 = 5'hc == index;
  assign T171 = ! T169;
  assign T172 = T174 ? 1'h0 : T173;
  assign T173 = Mapper_12_io_tx_val && Fifo_32_io_enq_rdy;
  assign T174 = ! T173;
  assign T175 = T178 ? 1'h0 : T176;
  assign T176 = T177 && Fifo_31_io_deq_val;
  assign T177 = 5'hb == index;
  assign T178 = ! T176;
  assign T179 = T181 ? 1'h0 : T180;
  assign T180 = Mapper_11_io_tx_val && Fifo_31_io_enq_rdy;
  assign T181 = ! T180;
  assign T182 = T185 ? 1'h0 : T183;
  assign T183 = T184 && Fifo_30_io_deq_val;
  assign T184 = 5'ha == index;
  assign T185 = ! T183;
  assign T186 = T188 ? 1'h0 : T187;
  assign T187 = Mapper_10_io_tx_val && Fifo_30_io_enq_rdy;
  assign T188 = ! T187;
  assign T189 = T192 ? 1'h0 : T190;
  assign T190 = T191 && Fifo_29_io_deq_val;
  assign T191 = 5'h9 == index;
  assign T192 = ! T190;
  assign T193 = T195 ? 1'h0 : T194;
  assign T194 = Mapper_9_io_tx_val && Fifo_29_io_enq_rdy;
  assign T195 = ! T194;
  assign T196 = T199 ? 1'h0 : T197;
  assign T197 = T198 && Fifo_28_io_deq_val;
  assign T198 = 5'h8 == index;
  assign T199 = ! T197;
  assign T200 = T202 ? 1'h0 : T201;
  assign T201 = Mapper_8_io_tx_val && Fifo_28_io_enq_rdy;
  assign T202 = ! T201;
  assign T203 = T206 ? 1'h0 : T204;
  assign T204 = T205 && Fifo_27_io_deq_val;
  assign T205 = 5'h7 == index;
  assign T206 = ! T204;
  assign T207 = T209 ? 1'h0 : T208;
  assign T208 = Mapper_7_io_tx_val && Fifo_27_io_enq_rdy;
  assign T209 = ! T208;
  assign T210 = T213 ? 1'h0 : T211;
  assign T211 = T212 && Fifo_26_io_deq_val;
  assign T212 = 5'h6 == index;
  assign T213 = ! T211;
  assign T214 = T216 ? 1'h0 : T215;
  assign T215 = Mapper_6_io_tx_val && Fifo_26_io_enq_rdy;
  assign T216 = ! T215;
  assign T217 = T220 ? 1'h0 : T218;
  assign T218 = T219 && Fifo_25_io_deq_val;
  assign T219 = 5'h5 == index;
  assign T220 = ! T218;
  assign T221 = T223 ? 1'h0 : T222;
  assign T222 = Mapper_5_io_tx_val && Fifo_25_io_enq_rdy;
  assign T223 = ! T222;
  assign T224 = T227 ? 1'h0 : T225;
  assign T225 = T226 && Fifo_24_io_deq_val;
  assign T226 = 5'h4 == index;
  assign T227 = ! T225;
  assign T228 = T230 ? 1'h0 : T229;
  assign T229 = Mapper_4_io_tx_val && Fifo_24_io_enq_rdy;
  assign T230 = ! T229;
  assign T231 = T234 ? 1'h0 : T232;
  assign T232 = T233 && Fifo_23_io_deq_val;
  assign T233 = 5'h3 == index;
  assign T234 = ! T232;
  assign T235 = T237 ? 1'h0 : T236;
  assign T236 = Mapper_3_io_tx_val && Fifo_23_io_enq_rdy;
  assign T237 = ! T236;
  assign T238 = T241 ? 1'h0 : T239;
  assign T239 = T240 && Fifo_22_io_deq_val;
  assign T240 = 5'h2 == index;
  assign T241 = ! T239;
  assign T242 = T244 ? 1'h0 : T243;
  assign T243 = Mapper_2_io_tx_val && Fifo_22_io_enq_rdy;
  assign T244 = ! T243;
  assign T245 = T248 ? 1'h0 : T246;
  assign T246 = T247 && Fifo_21_io_deq_val;
  assign T247 = 5'h1 == index;
  assign T248 = ! T246;
  assign T249 = T251 ? 1'h0 : T250;
  assign T250 = Mapper_1_io_tx_val && Fifo_21_io_enq_rdy;
  assign T251 = ! T250;
  assign T252 = T255 ? 1'h0 : T253;
  assign T253 = T254 && Fifo_20_io_deq_val;
  assign T254 = 5'h0 == index;
  assign T255 = ! T253;
  assign T256 = T258 ? 1'h0 : T257;
  assign T257 = Mapper_0_io_tx_val && Fifo_20_io_enq_rdy;
  assign T258 = ! T257;
  assign T259 = T2 ? 1'h0 : T1;
  assign T260 = T419 ? 1'h0 : T261;
  assign T261 = T262 && Fifo_19_io_enq_rdy;
  assign T262 = T263 && io_rx_val;
  assign T263 = 5'h13 == inCounter;
  assign T264 = T265 || T261;
  assign T265 = T269 || T266;
  assign T266 = T267 && Fifo_18_io_enq_rdy;
  assign T267 = T268 && io_rx_val;
  assign T268 = 5'h12 == inCounter;
  assign T269 = T273 || T270;
  assign T270 = T271 && Fifo_17_io_enq_rdy;
  assign T271 = T272 && io_rx_val;
  assign T272 = 5'h11 == inCounter;
  assign T273 = T277 || T274;
  assign T274 = T275 && Fifo_16_io_enq_rdy;
  assign T275 = T276 && io_rx_val;
  assign T276 = 5'h10 == inCounter;
  assign T277 = T281 || T278;
  assign T278 = T279 && Fifo_15_io_enq_rdy;
  assign T279 = T280 && io_rx_val;
  assign T280 = 5'hf == inCounter;
  assign T281 = T285 || T282;
  assign T282 = T283 && Fifo_14_io_enq_rdy;
  assign T283 = T284 && io_rx_val;
  assign T284 = 5'he == inCounter;
  assign T285 = T289 || T286;
  assign T286 = T287 && Fifo_13_io_enq_rdy;
  assign T287 = T288 && io_rx_val;
  assign T288 = 5'hd == inCounter;
  assign T289 = T293 || T290;
  assign T290 = T291 && Fifo_12_io_enq_rdy;
  assign T291 = T292 && io_rx_val;
  assign T292 = 5'hc == inCounter;
  assign T293 = T297 || T294;
  assign T294 = T295 && Fifo_11_io_enq_rdy;
  assign T295 = T296 && io_rx_val;
  assign T296 = 5'hb == inCounter;
  assign T297 = T301 || T298;
  assign T298 = T299 && Fifo_10_io_enq_rdy;
  assign T299 = T300 && io_rx_val;
  assign T300 = 5'ha == inCounter;
  assign T301 = T305 || T302;
  assign T302 = T303 && Fifo_9_io_enq_rdy;
  assign T303 = T304 && io_rx_val;
  assign T304 = 5'h9 == inCounter;
  assign T305 = T309 || T306;
  assign T306 = T307 && Fifo_8_io_enq_rdy;
  assign T307 = T308 && io_rx_val;
  assign T308 = 5'h8 == inCounter;
  assign T309 = T313 || T310;
  assign T310 = T311 && Fifo_7_io_enq_rdy;
  assign T311 = T312 && io_rx_val;
  assign T312 = 5'h7 == inCounter;
  assign T313 = T317 || T314;
  assign T314 = T315 && Fifo_6_io_enq_rdy;
  assign T315 = T316 && io_rx_val;
  assign T316 = 5'h6 == inCounter;
  assign T317 = T321 || T318;
  assign T318 = T319 && Fifo_5_io_enq_rdy;
  assign T319 = T320 && io_rx_val;
  assign T320 = 5'h5 == inCounter;
  assign T321 = T325 || T322;
  assign T322 = T323 && Fifo_4_io_enq_rdy;
  assign T323 = T324 && io_rx_val;
  assign T324 = 5'h4 == inCounter;
  assign T325 = T329 || T326;
  assign T326 = T327 && Fifo_3_io_enq_rdy;
  assign T327 = T328 && io_rx_val;
  assign T328 = 5'h3 == inCounter;
  assign T329 = T333 || T330;
  assign T330 = T331 && Fifo_2_io_enq_rdy;
  assign T331 = T332 && io_rx_val;
  assign T332 = 5'h2 == inCounter;
  assign T333 = T337 || T334;
  assign T334 = T335 && Fifo_1_io_enq_rdy;
  assign T335 = T336 && io_rx_val;
  assign T336 = 5'h1 == inCounter;
  assign T337 = T338 && Fifo_0_io_enq_rdy;
  assign T338 = T339 && io_rx_val;
  assign T339 = 5'h0 == inCounter;
  assign T340 = T261 ? T416 : T341;
  assign T341 = T266 ? T413 : T342;
  assign T342 = T270 ? T410 : T343;
  assign T343 = T274 ? T407 : T344;
  assign T344 = T278 ? T404 : T345;
  assign T345 = T282 ? T401 : T346;
  assign T346 = T286 ? T398 : T347;
  assign T347 = T290 ? T395 : T348;
  assign T348 = T294 ? T392 : T349;
  assign T349 = T298 ? T389 : T350;
  assign T350 = T302 ? T386 : T351;
  assign T351 = T306 ? T383 : T352;
  assign T352 = T310 ? T380 : T353;
  assign T353 = T314 ? T377 : T354;
  assign T354 = T318 ? T374 : T355;
  assign T355 = T322 ? T371 : T356;
  assign T356 = T326 ? T368 : T357;
  assign T357 = T330 ? T365 : T358;
  assign T358 = T334 ? T362 : T359;
  assign T359 = T361 ? 5'h0 : T360;
  assign T360 = inCounter + 5'h1;
  assign T361 = inCounter == 5'h13;
  assign T362 = T364 ? 5'h0 : T363;
  assign T363 = inCounter + 5'h1;
  assign T364 = inCounter == 5'h13;
  assign T365 = T367 ? 5'h0 : T366;
  assign T366 = inCounter + 5'h1;
  assign T367 = inCounter == 5'h13;
  assign T368 = T370 ? 5'h0 : T369;
  assign T369 = inCounter + 5'h1;
  assign T370 = inCounter == 5'h13;
  assign T371 = T373 ? 5'h0 : T372;
  assign T372 = inCounter + 5'h1;
  assign T373 = inCounter == 5'h13;
  assign T374 = T376 ? 5'h0 : T375;
  assign T375 = inCounter + 5'h1;
  assign T376 = inCounter == 5'h13;
  assign T377 = T379 ? 5'h0 : T378;
  assign T378 = inCounter + 5'h1;
  assign T379 = inCounter == 5'h13;
  assign T380 = T382 ? 5'h0 : T381;
  assign T381 = inCounter + 5'h1;
  assign T382 = inCounter == 5'h13;
  assign T383 = T385 ? 5'h0 : T384;
  assign T384 = inCounter + 5'h1;
  assign T385 = inCounter == 5'h13;
  assign T386 = T388 ? 5'h0 : T387;
  assign T387 = inCounter + 5'h1;
  assign T388 = inCounter == 5'h13;
  assign T389 = T391 ? 5'h0 : T390;
  assign T390 = inCounter + 5'h1;
  assign T391 = inCounter == 5'h13;
  assign T392 = T394 ? 5'h0 : T393;
  assign T393 = inCounter + 5'h1;
  assign T394 = inCounter == 5'h13;
  assign T395 = T397 ? 5'h0 : T396;
  assign T396 = inCounter + 5'h1;
  assign T397 = inCounter == 5'h13;
  assign T398 = T400 ? 5'h0 : T399;
  assign T399 = inCounter + 5'h1;
  assign T400 = inCounter == 5'h13;
  assign T401 = T403 ? 5'h0 : T402;
  assign T402 = inCounter + 5'h1;
  assign T403 = inCounter == 5'h13;
  assign T404 = T406 ? 5'h0 : T405;
  assign T405 = inCounter + 5'h1;
  assign T406 = inCounter == 5'h13;
  assign T407 = T409 ? 5'h0 : T408;
  assign T408 = inCounter + 5'h1;
  assign T409 = inCounter == 5'h13;
  assign T410 = T412 ? 5'h0 : T411;
  assign T411 = inCounter + 5'h1;
  assign T412 = inCounter == 5'h13;
  assign T413 = T415 ? 5'h0 : T414;
  assign T414 = inCounter + 5'h1;
  assign T415 = inCounter == 5'h13;
  assign T416 = T418 ? 5'h0 : T417;
  assign T417 = inCounter + 5'h1;
  assign T418 = inCounter == 5'h13;
  assign T419 = ! T261;
  assign T420 = T5 ? 1'h0 : T4;
  assign T421 = T422 ? 1'h0 : T266;
  assign T422 = ! T266;
  assign T423 = T8 ? 1'h0 : T7;
  assign T424 = T425 ? 1'h0 : T270;
  assign T425 = ! T270;
  assign T426 = T11 ? 1'h0 : T10;
  assign T427 = T428 ? 1'h0 : T274;
  assign T428 = ! T274;
  assign T429 = T14 ? 1'h0 : T13;
  assign T430 = T431 ? 1'h0 : T278;
  assign T431 = ! T278;
  assign T432 = T17 ? 1'h0 : T16;
  assign T433 = T434 ? 1'h0 : T282;
  assign T434 = ! T282;
  assign T435 = T20 ? 1'h0 : T19;
  assign T436 = T437 ? 1'h0 : T286;
  assign T437 = ! T286;
  assign T438 = T23 ? 1'h0 : T22;
  assign T439 = T440 ? 1'h0 : T290;
  assign T440 = ! T290;
  assign T441 = T26 ? 1'h0 : T25;
  assign T442 = T443 ? 1'h0 : T294;
  assign T443 = ! T294;
  assign T444 = T29 ? 1'h0 : T28;
  assign T445 = T446 ? 1'h0 : T298;
  assign T446 = ! T298;
  assign T447 = T32 ? 1'h0 : T31;
  assign T448 = T449 ? 1'h0 : T302;
  assign T449 = ! T302;
  assign T450 = T35 ? 1'h0 : T34;
  assign T451 = T452 ? 1'h0 : T306;
  assign T452 = ! T306;
  assign T453 = T38 ? 1'h0 : T37;
  assign T454 = T455 ? 1'h0 : T310;
  assign T455 = ! T310;
  assign T456 = T41 ? 1'h0 : T40;
  assign T457 = T458 ? 1'h0 : T314;
  assign T458 = ! T314;
  assign T459 = T44 ? 1'h0 : T43;
  assign T460 = T461 ? 1'h0 : T318;
  assign T461 = ! T318;
  assign T462 = T47 ? 1'h0 : T46;
  assign T463 = T464 ? 1'h0 : T322;
  assign T464 = ! T322;
  assign T465 = T50 ? 1'h0 : T49;
  assign T466 = T467 ? 1'h0 : T326;
  assign T467 = ! T326;
  assign T468 = T53 ? 1'h0 : T52;
  assign T469 = T470 ? 1'h0 : T330;
  assign T470 = ! T330;
  assign T471 = T56 ? 1'h0 : T55;
  assign T472 = T473 ? 1'h0 : T334;
  assign T473 = ! T334;
  assign T474 = T59 ? 1'h0 : T58;
  assign T475 = T476 ? 1'h0 : T337;
  assign T476 = ! T337;
  assign io_tx_val = T477;
  assign T477 = T61 ? 1'h1 : T478;
  assign T478 = T127 ? 1'h1 : T479;
  assign T479 = T134 ? 1'h1 : T480;
  assign T480 = T141 ? 1'h1 : T481;
  assign T481 = T148 ? 1'h1 : T482;
  assign T482 = T155 ? 1'h1 : T483;
  assign T483 = T162 ? 1'h1 : T484;
  assign T484 = T169 ? 1'h1 : T485;
  assign T485 = T176 ? 1'h1 : T486;
  assign T486 = T183 ? 1'h1 : T487;
  assign T487 = T190 ? 1'h1 : T488;
  assign T488 = T197 ? 1'h1 : T489;
  assign T489 = T204 ? 1'h1 : T490;
  assign T490 = T211 ? 1'h1 : T491;
  assign T491 = T218 ? 1'h1 : T492;
  assign T492 = T225 ? 1'h1 : T493;
  assign T493 = T232 ? 1'h1 : T494;
  assign T494 = T239 ? 1'h1 : T495;
  assign T495 = T246 ? 1'h1 : T253;
  assign io_tx_dat_int = T496;
  assign T496 = T61 ? Fifo_39_io_deq_dat_int : T497;
  assign T497 = T127 ? Fifo_38_io_deq_dat_int : T498;
  assign T498 = T134 ? Fifo_37_io_deq_dat_int : T499;
  assign T499 = T141 ? Fifo_36_io_deq_dat_int : T500;
  assign T500 = T148 ? Fifo_35_io_deq_dat_int : T501;
  assign T501 = T155 ? Fifo_34_io_deq_dat_int : T502;
  assign T502 = T162 ? Fifo_33_io_deq_dat_int : T503;
  assign T503 = T169 ? Fifo_32_io_deq_dat_int : T504;
  assign T504 = T176 ? Fifo_31_io_deq_dat_int : T505;
  assign T505 = T183 ? Fifo_30_io_deq_dat_int : T506;
  assign T506 = T190 ? Fifo_29_io_deq_dat_int : T507;
  assign T507 = T197 ? Fifo_28_io_deq_dat_int : T508;
  assign T508 = T204 ? Fifo_27_io_deq_dat_int : T509;
  assign T509 = T211 ? Fifo_26_io_deq_dat_int : T510;
  assign T510 = T218 ? Fifo_25_io_deq_dat_int : T511;
  assign T511 = T225 ? Fifo_24_io_deq_dat_int : T512;
  assign T512 = T232 ? Fifo_23_io_deq_dat_int : T513;
  assign T513 = T239 ? Fifo_22_io_deq_dat_int : T514;
  assign T514 = T246 ? Fifo_21_io_deq_dat_int : T515;
  assign T515 = T253 ? Fifo_20_io_deq_dat_int : 64'h0;
  Fifo_1 Fifo_0(.clk(clk), .reset(reset),
       .io_enq_val( T475 ),
       .io_enq_rdy( Fifo_0_io_enq_rdy ),
       .io_deq_val( Fifo_0_io_deq_val ),
       .io_deq_rdy( T474 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_0_io_deq_dat_int )
  );
  Fifo_1 Fifo_1(.clk(clk), .reset(reset),
       .io_enq_val( T472 ),
       .io_enq_rdy( Fifo_1_io_enq_rdy ),
       .io_deq_val( Fifo_1_io_deq_val ),
       .io_deq_rdy( T471 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_1_io_deq_dat_int )
  );
  Fifo_1 Fifo_2(.clk(clk), .reset(reset),
       .io_enq_val( T469 ),
       .io_enq_rdy( Fifo_2_io_enq_rdy ),
       .io_deq_val( Fifo_2_io_deq_val ),
       .io_deq_rdy( T468 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_2_io_deq_dat_int )
  );
  Fifo_1 Fifo_3(.clk(clk), .reset(reset),
       .io_enq_val( T466 ),
       .io_enq_rdy( Fifo_3_io_enq_rdy ),
       .io_deq_val( Fifo_3_io_deq_val ),
       .io_deq_rdy( T465 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_3_io_deq_dat_int )
  );
  Fifo_1 Fifo_4(.clk(clk), .reset(reset),
       .io_enq_val( T463 ),
       .io_enq_rdy( Fifo_4_io_enq_rdy ),
       .io_deq_val( Fifo_4_io_deq_val ),
       .io_deq_rdy( T462 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_4_io_deq_dat_int )
  );
  Fifo_1 Fifo_5(.clk(clk), .reset(reset),
       .io_enq_val( T460 ),
       .io_enq_rdy( Fifo_5_io_enq_rdy ),
       .io_deq_val( Fifo_5_io_deq_val ),
       .io_deq_rdy( T459 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_5_io_deq_dat_int )
  );
  Fifo_1 Fifo_6(.clk(clk), .reset(reset),
       .io_enq_val( T457 ),
       .io_enq_rdy( Fifo_6_io_enq_rdy ),
       .io_deq_val( Fifo_6_io_deq_val ),
       .io_deq_rdy( T456 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_6_io_deq_dat_int )
  );
  Fifo_1 Fifo_7(.clk(clk), .reset(reset),
       .io_enq_val( T454 ),
       .io_enq_rdy( Fifo_7_io_enq_rdy ),
       .io_deq_val( Fifo_7_io_deq_val ),
       .io_deq_rdy( T453 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_7_io_deq_dat_int )
  );
  Fifo_1 Fifo_8(.clk(clk), .reset(reset),
       .io_enq_val( T451 ),
       .io_enq_rdy( Fifo_8_io_enq_rdy ),
       .io_deq_val( Fifo_8_io_deq_val ),
       .io_deq_rdy( T450 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_8_io_deq_dat_int )
  );
  Fifo_1 Fifo_9(.clk(clk), .reset(reset),
       .io_enq_val( T448 ),
       .io_enq_rdy( Fifo_9_io_enq_rdy ),
       .io_deq_val( Fifo_9_io_deq_val ),
       .io_deq_rdy( T447 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_9_io_deq_dat_int )
  );
  Fifo_1 Fifo_10(.clk(clk), .reset(reset),
       .io_enq_val( T445 ),
       .io_enq_rdy( Fifo_10_io_enq_rdy ),
       .io_deq_val( Fifo_10_io_deq_val ),
       .io_deq_rdy( T444 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_10_io_deq_dat_int )
  );
  Fifo_1 Fifo_11(.clk(clk), .reset(reset),
       .io_enq_val( T442 ),
       .io_enq_rdy( Fifo_11_io_enq_rdy ),
       .io_deq_val( Fifo_11_io_deq_val ),
       .io_deq_rdy( T441 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_11_io_deq_dat_int )
  );
  Fifo_1 Fifo_12(.clk(clk), .reset(reset),
       .io_enq_val( T439 ),
       .io_enq_rdy( Fifo_12_io_enq_rdy ),
       .io_deq_val( Fifo_12_io_deq_val ),
       .io_deq_rdy( T438 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_12_io_deq_dat_int )
  );
  Fifo_1 Fifo_13(.clk(clk), .reset(reset),
       .io_enq_val( T436 ),
       .io_enq_rdy( Fifo_13_io_enq_rdy ),
       .io_deq_val( Fifo_13_io_deq_val ),
       .io_deq_rdy( T435 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_13_io_deq_dat_int )
  );
  Fifo_1 Fifo_14(.clk(clk), .reset(reset),
       .io_enq_val( T433 ),
       .io_enq_rdy( Fifo_14_io_enq_rdy ),
       .io_deq_val( Fifo_14_io_deq_val ),
       .io_deq_rdy( T432 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_14_io_deq_dat_int )
  );
  Fifo_1 Fifo_15(.clk(clk), .reset(reset),
       .io_enq_val( T430 ),
       .io_enq_rdy( Fifo_15_io_enq_rdy ),
       .io_deq_val( Fifo_15_io_deq_val ),
       .io_deq_rdy( T429 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_15_io_deq_dat_int )
  );
  Fifo_1 Fifo_16(.clk(clk), .reset(reset),
       .io_enq_val( T427 ),
       .io_enq_rdy( Fifo_16_io_enq_rdy ),
       .io_deq_val( Fifo_16_io_deq_val ),
       .io_deq_rdy( T426 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_16_io_deq_dat_int )
  );
  Fifo_1 Fifo_17(.clk(clk), .reset(reset),
       .io_enq_val( T424 ),
       .io_enq_rdy( Fifo_17_io_enq_rdy ),
       .io_deq_val( Fifo_17_io_deq_val ),
       .io_deq_rdy( T423 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_17_io_deq_dat_int )
  );
  Fifo_1 Fifo_18(.clk(clk), .reset(reset),
       .io_enq_val( T421 ),
       .io_enq_rdy( Fifo_18_io_enq_rdy ),
       .io_deq_val( Fifo_18_io_deq_val ),
       .io_deq_rdy( T420 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_18_io_deq_dat_int )
  );
  Fifo_1 Fifo_19(.clk(clk), .reset(reset),
       .io_enq_val( T260 ),
       .io_enq_rdy( Fifo_19_io_enq_rdy ),
       .io_deq_val( Fifo_19_io_deq_val ),
       .io_deq_rdy( T259 ),
       .io_enq_dat_int( io_rx_dat_int ),
       .io_deq_dat_int( Fifo_19_io_deq_dat_int )
  );
  Fifo_1 Fifo_20(.clk(clk), .reset(reset),
       .io_enq_val( T256 ),
       .io_enq_rdy( Fifo_20_io_enq_rdy ),
       .io_deq_val( Fifo_20_io_deq_val ),
       .io_deq_rdy( T252 ),
       .io_enq_dat_int( Mapper_0_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_20_io_deq_dat_int )
  );
  Fifo_1 Fifo_21(.clk(clk), .reset(reset),
       .io_enq_val( T249 ),
       .io_enq_rdy( Fifo_21_io_enq_rdy ),
       .io_deq_val( Fifo_21_io_deq_val ),
       .io_deq_rdy( T245 ),
       .io_enq_dat_int( Mapper_1_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_21_io_deq_dat_int )
  );
  Fifo_1 Fifo_22(.clk(clk), .reset(reset),
       .io_enq_val( T242 ),
       .io_enq_rdy( Fifo_22_io_enq_rdy ),
       .io_deq_val( Fifo_22_io_deq_val ),
       .io_deq_rdy( T238 ),
       .io_enq_dat_int( Mapper_2_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_22_io_deq_dat_int )
  );
  Fifo_1 Fifo_23(.clk(clk), .reset(reset),
       .io_enq_val( T235 ),
       .io_enq_rdy( Fifo_23_io_enq_rdy ),
       .io_deq_val( Fifo_23_io_deq_val ),
       .io_deq_rdy( T231 ),
       .io_enq_dat_int( Mapper_3_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_23_io_deq_dat_int )
  );
  Fifo_1 Fifo_24(.clk(clk), .reset(reset),
       .io_enq_val( T228 ),
       .io_enq_rdy( Fifo_24_io_enq_rdy ),
       .io_deq_val( Fifo_24_io_deq_val ),
       .io_deq_rdy( T224 ),
       .io_enq_dat_int( Mapper_4_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_24_io_deq_dat_int )
  );
  Fifo_1 Fifo_25(.clk(clk), .reset(reset),
       .io_enq_val( T221 ),
       .io_enq_rdy( Fifo_25_io_enq_rdy ),
       .io_deq_val( Fifo_25_io_deq_val ),
       .io_deq_rdy( T217 ),
       .io_enq_dat_int( Mapper_5_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_25_io_deq_dat_int )
  );
  Fifo_1 Fifo_26(.clk(clk), .reset(reset),
       .io_enq_val( T214 ),
       .io_enq_rdy( Fifo_26_io_enq_rdy ),
       .io_deq_val( Fifo_26_io_deq_val ),
       .io_deq_rdy( T210 ),
       .io_enq_dat_int( Mapper_6_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_26_io_deq_dat_int )
  );
  Fifo_1 Fifo_27(.clk(clk), .reset(reset),
       .io_enq_val( T207 ),
       .io_enq_rdy( Fifo_27_io_enq_rdy ),
       .io_deq_val( Fifo_27_io_deq_val ),
       .io_deq_rdy( T203 ),
       .io_enq_dat_int( Mapper_7_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_27_io_deq_dat_int )
  );
  Fifo_1 Fifo_28(.clk(clk), .reset(reset),
       .io_enq_val( T200 ),
       .io_enq_rdy( Fifo_28_io_enq_rdy ),
       .io_deq_val( Fifo_28_io_deq_val ),
       .io_deq_rdy( T196 ),
       .io_enq_dat_int( Mapper_8_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_28_io_deq_dat_int )
  );
  Fifo_1 Fifo_29(.clk(clk), .reset(reset),
       .io_enq_val( T193 ),
       .io_enq_rdy( Fifo_29_io_enq_rdy ),
       .io_deq_val( Fifo_29_io_deq_val ),
       .io_deq_rdy( T189 ),
       .io_enq_dat_int( Mapper_9_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_29_io_deq_dat_int )
  );
  Fifo_1 Fifo_30(.clk(clk), .reset(reset),
       .io_enq_val( T186 ),
       .io_enq_rdy( Fifo_30_io_enq_rdy ),
       .io_deq_val( Fifo_30_io_deq_val ),
       .io_deq_rdy( T182 ),
       .io_enq_dat_int( Mapper_10_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_30_io_deq_dat_int )
  );
  Fifo_1 Fifo_31(.clk(clk), .reset(reset),
       .io_enq_val( T179 ),
       .io_enq_rdy( Fifo_31_io_enq_rdy ),
       .io_deq_val( Fifo_31_io_deq_val ),
       .io_deq_rdy( T175 ),
       .io_enq_dat_int( Mapper_11_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_31_io_deq_dat_int )
  );
  Fifo_1 Fifo_32(.clk(clk), .reset(reset),
       .io_enq_val( T172 ),
       .io_enq_rdy( Fifo_32_io_enq_rdy ),
       .io_deq_val( Fifo_32_io_deq_val ),
       .io_deq_rdy( T168 ),
       .io_enq_dat_int( Mapper_12_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_32_io_deq_dat_int )
  );
  Fifo_1 Fifo_33(.clk(clk), .reset(reset),
       .io_enq_val( T165 ),
       .io_enq_rdy( Fifo_33_io_enq_rdy ),
       .io_deq_val( Fifo_33_io_deq_val ),
       .io_deq_rdy( T161 ),
       .io_enq_dat_int( Mapper_13_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_33_io_deq_dat_int )
  );
  Fifo_1 Fifo_34(.clk(clk), .reset(reset),
       .io_enq_val( T158 ),
       .io_enq_rdy( Fifo_34_io_enq_rdy ),
       .io_deq_val( Fifo_34_io_deq_val ),
       .io_deq_rdy( T154 ),
       .io_enq_dat_int( Mapper_14_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_34_io_deq_dat_int )
  );
  Fifo_1 Fifo_35(.clk(clk), .reset(reset),
       .io_enq_val( T151 ),
       .io_enq_rdy( Fifo_35_io_enq_rdy ),
       .io_deq_val( Fifo_35_io_deq_val ),
       .io_deq_rdy( T147 ),
       .io_enq_dat_int( Mapper_15_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_35_io_deq_dat_int )
  );
  Fifo_1 Fifo_36(.clk(clk), .reset(reset),
       .io_enq_val( T144 ),
       .io_enq_rdy( Fifo_36_io_enq_rdy ),
       .io_deq_val( Fifo_36_io_deq_val ),
       .io_deq_rdy( T140 ),
       .io_enq_dat_int( Mapper_16_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_36_io_deq_dat_int )
  );
  Fifo_1 Fifo_37(.clk(clk), .reset(reset),
       .io_enq_val( T137 ),
       .io_enq_rdy( Fifo_37_io_enq_rdy ),
       .io_deq_val( Fifo_37_io_deq_val ),
       .io_deq_rdy( T133 ),
       .io_enq_dat_int( Mapper_17_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_37_io_deq_dat_int )
  );
  Fifo_1 Fifo_38(.clk(clk), .reset(reset),
       .io_enq_val( T130 ),
       .io_enq_rdy( Fifo_38_io_enq_rdy ),
       .io_deq_val( Fifo_38_io_deq_val ),
       .io_deq_rdy( T126 ),
       .io_enq_dat_int( Mapper_18_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_38_io_deq_dat_int )
  );
  Fifo_1 Fifo_39(.clk(clk), .reset(reset),
       .io_enq_val( T123 ),
       .io_enq_rdy( Fifo_39_io_enq_rdy ),
       .io_deq_val( Fifo_39_io_deq_val ),
       .io_deq_rdy( T60 ),
       .io_enq_dat_int( Mapper_19_io_tx_dat_int ),
       .io_deq_dat_int( Fifo_39_io_deq_dat_int )
  );
  Mapper Mapper_0(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_0_io_deq_dat_int ),
       .io_rx_val( T57 ),
       .io_rx_rdy( Mapper_0_io_rx_rdy ),
       .io_tx_dat_int( Mapper_0_io_tx_dat_int ),
       .io_tx_val( Mapper_0_io_tx_val )
  );
  Mapper Mapper_1(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_1_io_deq_dat_int ),
       .io_rx_val( T54 ),
       .io_rx_rdy( Mapper_1_io_rx_rdy ),
       .io_tx_dat_int( Mapper_1_io_tx_dat_int ),
       .io_tx_val( Mapper_1_io_tx_val )
  );
  Mapper Mapper_2(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_2_io_deq_dat_int ),
       .io_rx_val( T51 ),
       .io_rx_rdy( Mapper_2_io_rx_rdy ),
       .io_tx_dat_int( Mapper_2_io_tx_dat_int ),
       .io_tx_val( Mapper_2_io_tx_val )
  );
  Mapper Mapper_3(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_3_io_deq_dat_int ),
       .io_rx_val( T48 ),
       .io_rx_rdy( Mapper_3_io_rx_rdy ),
       .io_tx_dat_int( Mapper_3_io_tx_dat_int ),
       .io_tx_val( Mapper_3_io_tx_val )
  );
  Mapper Mapper_4(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_4_io_deq_dat_int ),
       .io_rx_val( T45 ),
       .io_rx_rdy( Mapper_4_io_rx_rdy ),
       .io_tx_dat_int( Mapper_4_io_tx_dat_int ),
       .io_tx_val( Mapper_4_io_tx_val )
  );
  Mapper Mapper_5(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_5_io_deq_dat_int ),
       .io_rx_val( T42 ),
       .io_rx_rdy( Mapper_5_io_rx_rdy ),
       .io_tx_dat_int( Mapper_5_io_tx_dat_int ),
       .io_tx_val( Mapper_5_io_tx_val )
  );
  Mapper Mapper_6(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_6_io_deq_dat_int ),
       .io_rx_val( T39 ),
       .io_rx_rdy( Mapper_6_io_rx_rdy ),
       .io_tx_dat_int( Mapper_6_io_tx_dat_int ),
       .io_tx_val( Mapper_6_io_tx_val )
  );
  Mapper Mapper_7(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_7_io_deq_dat_int ),
       .io_rx_val( T36 ),
       .io_rx_rdy( Mapper_7_io_rx_rdy ),
       .io_tx_dat_int( Mapper_7_io_tx_dat_int ),
       .io_tx_val( Mapper_7_io_tx_val )
  );
  Mapper Mapper_8(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_8_io_deq_dat_int ),
       .io_rx_val( T33 ),
       .io_rx_rdy( Mapper_8_io_rx_rdy ),
       .io_tx_dat_int( Mapper_8_io_tx_dat_int ),
       .io_tx_val( Mapper_8_io_tx_val )
  );
  Mapper Mapper_9(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_9_io_deq_dat_int ),
       .io_rx_val( T30 ),
       .io_rx_rdy( Mapper_9_io_rx_rdy ),
       .io_tx_dat_int( Mapper_9_io_tx_dat_int ),
       .io_tx_val( Mapper_9_io_tx_val )
  );
  Mapper Mapper_10(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_10_io_deq_dat_int ),
       .io_rx_val( T27 ),
       .io_rx_rdy( Mapper_10_io_rx_rdy ),
       .io_tx_dat_int( Mapper_10_io_tx_dat_int ),
       .io_tx_val( Mapper_10_io_tx_val )
  );
  Mapper Mapper_11(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_11_io_deq_dat_int ),
       .io_rx_val( T24 ),
       .io_rx_rdy( Mapper_11_io_rx_rdy ),
       .io_tx_dat_int( Mapper_11_io_tx_dat_int ),
       .io_tx_val( Mapper_11_io_tx_val )
  );
  Mapper Mapper_12(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_12_io_deq_dat_int ),
       .io_rx_val( T21 ),
       .io_rx_rdy( Mapper_12_io_rx_rdy ),
       .io_tx_dat_int( Mapper_12_io_tx_dat_int ),
       .io_tx_val( Mapper_12_io_tx_val )
  );
  Mapper Mapper_13(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_13_io_deq_dat_int ),
       .io_rx_val( T18 ),
       .io_rx_rdy( Mapper_13_io_rx_rdy ),
       .io_tx_dat_int( Mapper_13_io_tx_dat_int ),
       .io_tx_val( Mapper_13_io_tx_val )
  );
  Mapper Mapper_14(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_14_io_deq_dat_int ),
       .io_rx_val( T15 ),
       .io_rx_rdy( Mapper_14_io_rx_rdy ),
       .io_tx_dat_int( Mapper_14_io_tx_dat_int ),
       .io_tx_val( Mapper_14_io_tx_val )
  );
  Mapper Mapper_15(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_15_io_deq_dat_int ),
       .io_rx_val( T12 ),
       .io_rx_rdy( Mapper_15_io_rx_rdy ),
       .io_tx_dat_int( Mapper_15_io_tx_dat_int ),
       .io_tx_val( Mapper_15_io_tx_val )
  );
  Mapper Mapper_16(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_16_io_deq_dat_int ),
       .io_rx_val( T9 ),
       .io_rx_rdy( Mapper_16_io_rx_rdy ),
       .io_tx_dat_int( Mapper_16_io_tx_dat_int ),
       .io_tx_val( Mapper_16_io_tx_val )
  );
  Mapper Mapper_17(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_17_io_deq_dat_int ),
       .io_rx_val( T6 ),
       .io_rx_rdy( Mapper_17_io_rx_rdy ),
       .io_tx_dat_int( Mapper_17_io_tx_dat_int ),
       .io_tx_val( Mapper_17_io_tx_val )
  );
  Mapper Mapper_18(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_18_io_deq_dat_int ),
       .io_rx_val( T3 ),
       .io_rx_rdy( Mapper_18_io_rx_rdy ),
       .io_tx_dat_int( Mapper_18_io_tx_dat_int ),
       .io_tx_val( Mapper_18_io_tx_val )
  );
  Mapper Mapper_19(.clk(clk), .reset(reset),
       .io_rx_dat_int( Fifo_19_io_deq_dat_int ),
       .io_rx_val( T0 ),
       .io_rx_rdy( Mapper_19_io_rx_rdy ),
       .io_tx_dat_int( Mapper_19_io_tx_dat_int ),
       .io_tx_val( Mapper_19_io_tx_val )
  );

  always @(posedge clk) begin
    if(reset) begin
      inCounter <= 5'h0;
    end else if(T264) begin
      inCounter <= T340;
    end
  end
endmodule

module MrSimSimulation(input clk, input reset,
    input [63:0] io_enq_dat,
    input  io_enq_val,
    output io_enq_rdy,
    output[63:0] io_deq_dat,
    output io_deq_val,
    input  io_deq_rdy
);

  wire decode_io_tx_val;
  wire[63:0] decode_io_tx_dat_int;
  wire T0;
  wire decode_io_rx_rdy;
  wire Fifo_0_io_deq_val;
  wire[63:0] Fifo_0_io_deq_dat;
  wire Controller_io_tx_val;
  wire[63:0] Controller_io_tx_dat_int;
  wire[63:0] encode_io_tx_dat;
  wire encode_io_tx_val;
  wire T1;
  wire Fifo_1_io_deq_val;
  wire[63:0] Fifo_1_io_deq_dat;
  wire Fifo_0_io_enq_rdy;

  assign T0 = Fifo_0_io_deq_val && decode_io_rx_rdy;
  assign T1 = decode_io_rx_rdy && Fifo_0_io_deq_val;
  assign io_deq_val = Fifo_1_io_deq_val;
  assign io_deq_dat = Fifo_1_io_deq_dat;
  assign io_enq_rdy = Fifo_0_io_enq_rdy;
  Fifo_0 Fifo_0(.clk(clk), .reset(reset),
       .io_enq_val( io_enq_val ),
       .io_enq_rdy( Fifo_0_io_enq_rdy ),
       .io_deq_val( Fifo_0_io_deq_val ),
       .io_deq_rdy( T1 ),
       .io_enq_dat( io_enq_dat ),
       .io_deq_dat( Fifo_0_io_deq_dat )
  );
  Fifo_0 Fifo_1(.clk(clk), .reset(reset),
       .io_enq_val( encode_io_tx_val ),
       //.io_enq_rdy(  )
       .io_deq_val( Fifo_1_io_deq_val ),
       .io_deq_rdy( io_deq_rdy ),
       .io_enq_dat( encode_io_tx_dat ),
       .io_deq_dat( Fifo_1_io_deq_dat )
  );
  encode encode(
       .io_rx_dat_int( Controller_io_tx_dat_int ),
       //.io_rx_rdy(  )
       .io_rx_val( Controller_io_tx_val ),
       .io_tx_dat( encode_io_tx_dat ),
       .io_tx_val( encode_io_tx_val )
  );
  decode decode(
       .io_rx_dat( Fifo_0_io_deq_dat ),
       .io_rx_rdy( decode_io_rx_rdy ),
       .io_rx_val( T0 ),
       .io_tx_dat_int( decode_io_tx_dat_int ),
       .io_tx_val( decode_io_tx_val )
  );
  Controller Controller(.clk(clk), .reset(reset),
       .io_rx_dat_int( decode_io_tx_dat_int ),
       .io_rx_val( decode_io_tx_val ),
       .io_tx_dat_int( Controller_io_tx_dat_int ),
       .io_tx_val( Controller_io_tx_val )
  );
endmodule

